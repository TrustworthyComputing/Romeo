module s1423(VDD,CK,G0,G1,G10,G11,G12,G13,G14,G15,G16,G2,G3,G4,G5,G6,G7,
  G701BF,G702,G726,G727,G729,G8,G9);
input VDD,CK,G0,G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16;
output G726,G729,G702,G727,G701BF;

  wire G22,G332BF,G23,G328BF,G24,G109,G25,G113,G26,G118,G27,G125,G28,G129,G29,
    G140,G30,G144,G31,G149,G32,G154,G33,G159,G34,G166,G35,G175,G36,G189,G37,
    G193,G38,G198,G39,G208,G40,G214,G41,G218,G42,G237,G43,G242,G44,G247,G45,
    G252,G46,G260,G47,G303,G48,G309,G49,G315,G50,G321,G51,G360,G52,G365,G53,
    G373,G54,G379,G55,G384,G56,G392,G57,G397,G58,G405,G59,G408,G60,G416,G61,
    G424,G62,G427,G63,G438,G64,G441,G65,G447,G66,G451,G67,G459,G68,G464,G69,
    G469,G70,G477,G71,G494,G72,G498,G73,G503,G74,G526,G75,G531,G76,G536,G77,
    G541,G78,G548,G79,G565,G80,G569,G81,G573,G82,G577,G83,G590,G84,G608,G85,
    G613,G86,G657,G87,G663,G88,G669,G89,G675,G90,G682,G91,G687,G92,G693,G93,
    G705,G94,G707,G95,G713,II1,G332,II12,G328,G108,G712,G111,G112,G117,G124,
    G127,G128,G139,G142,G143,G148,G153,G158,G165,G174,G176,G178,G179,G180,G188,
    G191,G192,G197,G204,G207,G210,G213,G216,G217,G236,G259,G241,G246,G251,G258,
    G296,G297,G302,G305,G324,G308,G311,G314,G317,G320,G323,G336,G355,G339,G343,
    G348,G347,G351,G645,G354,G359,G372,G364,G371,G378,G391,G383,G390,G396,G404,
    G403,G407,G415,G423,G422,G426,G437,G440,G445,G446,G449,G450,G455,G456,G458,
    G476,G463,G468,G475,G486,G491,G500,G495,G499,G504,G511,G507,G510,G525,G589,
    G530,G535,G540,G547,G562,G610,G566,G570,G574,G588,G595,G593,G596,G597,G600,
    G601,G605,G609,G614,G615,G616,G617,G620,G623,G626,G629,G632,G635,G638,G641,
    G644,G656,G658,G659,II1162,G661,G662,G665,G678,G668,G671,G674,G677,II1183,
    G685,G696,G689,G695,II1203,G701,II1211,G704,G706,G711,G714,II1227,G715,
    II1230,G716,II1233,G717,II1236,G718,II1239,G719,II1242,G720,II1245,G721,
    II1248,G722,II1251,G723,II1254,G724,II1257,G725,II1260,II1264,G728,II1267,
    G101,G630,G631,G102,G633,G634,G103,G636,G637,G104,G639,G640,G105,G642,G643,
    G106,G114,G116,G133,G119,G121,G134,G122,G130,G132,G136,G700,G135,G137,G145,
    G147,G168,G150,G152,G169,G155,G157,G170,G160,G162,G171,G163,G177,G172,G173,
    G185,G181,G182,G186,G194,G196,G202,G199,G201,G203,G522,G205,G211,G219,G221,
    G223,G222,G183,G224,G225,G226,G227,G228,G229,G432,G238,G240,G299,G243,G245,
    G262,G248,G250,G263,G253,G255,G264,G624,G625,G256,G261,G265,G271,G275,G266,
    G272,G276,G277,G273,G278,G279,G274,G280,G281,G304,G306,G307,G310,G312,G313,
    G316,G318,G319,G322,G325,G326,G329,G331,G330,G335,G337,G338,G342,G344,G345,
    G346,G349,G350,G358,G523,G361,G363,G366,G368,G375,G369,G374,G376,G377,G380,
    G382,G385,G387,G394,G388,G393,G395,G398,G400,G401,G406,G412,G409,G411,G413,
    G414,G417,G419,G420,G425,G431,G428,G430,G433,G356,G357,G435,G340,G341,G436,
    G352,G353,G439,G442,G443,G448,G452,G453,G457,G460,G462,G434,G465,G467,G479,
    G470,G472,G480,G473,G478,G481,G488,G505,G506,G489,G508,G509,G490,G512,G513,
    G492,G493,G496,G497,G501,G502,G527,G529,G604,G532,G534,G550,G537,G539,G551,
    G542,G544,G552,G545,G549,G553,G563,G564,G567,G568,G571,G572,G575,G576,G627,
    G628,G591,G592,G594,G621,G622,G524,G606,G607,G611,G612,G648,G646,G647,G649,
    G618,G619,G650,G651,G652,G653,G654,G655,G664,G666,G667,G670,G672,G673,G676,
    G679,G680,G683,G684,G688,G690,G691,G694,G697,G698,G703,G230,G708,G709,G599,
    G110,G126,G141,G167,G184,G190,G209,G215,G235,G233,G267,G268,G269,G282,G283,
    G270,G291,G292,G293,G294,G295,G300,G333,G334,G301,G518,G519,G520,G521,G487,
    G554,G555,G583,G584,G585,G586,G587,G561,G602,G603,G96,G97,G98,G99,G100,
    G681,G699,G686,G692,G107,G123,G138,G164,G187,G206,G212,G234,G231,G232,G298,
    G286,G287,G288,G284,G285,G289,G290,G482,G514,G483,G515,G484,G516,G485,G517,
    G556,G557,G558,G559,G560,G578,G579,G580,G581,G582,G598,G115,G120,G131,G146,
    G151,G156,G161,G195,G200,G220,G239,G244,G249,G254,G257,G327,G362,G367,G370,
    G381,G386,G389,G399,G402,G410,G418,G421,G429,G444,G454,G461,G466,G471,G474,
    G528,G533,G538,G543,G546,G660,G710;

  FD1 DFF_0(CK,G22,G332BF);
  FD1 DFF_1(CK,G23,G328BF);
  FD1 DFF_2(CK,G24,G109);
  FD1 DFF_3(CK,G25,G113);
  FD1 DFF_4(CK,G26,G118);
  FD1 DFF_5(CK,G27,G125);
  FD1 DFF_6(CK,G28,G129);
  FD1 DFF_7(CK,G29,G140);
  FD1 DFF_8(CK,G30,G144);
  FD1 DFF_9(CK,G31,G149);
  FD1 DFF_10(CK,G32,G154);
  FD1 DFF_11(CK,G33,G159);
  FD1 DFF_12(CK,G34,G166);
  FD1 DFF_13(CK,G35,G175);
  FD1 DFF_14(CK,G36,G189);
  FD1 DFF_15(CK,G37,G193);
  FD1 DFF_16(CK,G38,G198);
  FD1 DFF_17(CK,G39,G208);
  FD1 DFF_18(CK,G40,G214);
  FD1 DFF_19(CK,G41,G218);
  FD1 DFF_20(CK,G42,G237);
  FD1 DFF_21(CK,G43,G242);
  FD1 DFF_22(CK,G44,G247);
  FD1 DFF_23(CK,G45,G252);
  FD1 DFF_24(CK,G46,G260);
  FD1 DFF_25(CK,G47,G303);
  FD1 DFF_26(CK,G48,G309);
  FD1 DFF_27(CK,G49,G315);
  FD1 DFF_28(CK,G50,G321);
  FD1 DFF_29(CK,G51,G360);
  FD1 DFF_30(CK,G52,G365);
  FD1 DFF_31(CK,G53,G373);
  FD1 DFF_32(CK,G54,G379);
  FD1 DFF_33(CK,G55,G384);
  FD1 DFF_34(CK,G56,G392);
  FD1 DFF_35(CK,G57,G397);
  FD1 DFF_36(CK,G58,G405);
  FD1 DFF_37(CK,G59,G408);
  FD1 DFF_38(CK,G60,G416);
  FD1 DFF_39(CK,G61,G424);
  FD1 DFF_40(CK,G62,G427);
  FD1 DFF_41(CK,G63,G438);
  FD1 DFF_42(CK,G64,G441);
  FD1 DFF_43(CK,G65,G447);
  FD1 DFF_44(CK,G66,G451);
  FD1 DFF_45(CK,G67,G459);
  FD1 DFF_46(CK,G68,G464);
  FD1 DFF_47(CK,G69,G469);
  FD1 DFF_48(CK,G70,G477);
  FD1 DFF_49(CK,G71,G494);
  FD1 DFF_50(CK,G72,G498);
  FD1 DFF_51(CK,G73,G503);
  FD1 DFF_52(CK,G74,G526);
  FD1 DFF_53(CK,G75,G531);
  FD1 DFF_54(CK,G76,G536);
  FD1 DFF_55(CK,G77,G541);
  FD1 DFF_56(CK,G78,G548);
  FD1 DFF_57(CK,G79,G565);
  FD1 DFF_58(CK,G80,G569);
  FD1 DFF_59(CK,G81,G573);
  FD1 DFF_60(CK,G82,G577);
  FD1 DFF_61(CK,G83,G590);
  FD1 DFF_62(CK,G84,G608);
  FD1 DFF_63(CK,G85,G613);
  FD1 DFF_64(CK,G86,G657);
  FD1 DFF_65(CK,G87,G663);
  FD1 DFF_66(CK,G88,G669);
  FD1 DFF_67(CK,G89,G675);
  FD1 DFF_68(CK,G90,G682);
  FD1 DFF_69(CK,G91,G687);
  FD1 DFF_70(CK,G92,G693);
  FD1 DFF_71(CK,G93,G705);
  FD1 DFF_72(CK,G94,G707);
  FD1 DFF_73(CK,G95,G713);
  IV  NOT_0(II1,G332);
  IV  NOT_1(G332BF,II1);
  IV  NOT_2(II12,G328);
  IV  NOT_3(G328BF,II12);
  IV  NOT_4(G108,G712);
  IV  NOT_5(G111,G24);
  IV  NOT_6(G112,G712);
  IV  NOT_7(G117,G712);
  IV  NOT_8(G124,G712);
  IV  NOT_9(G127,G27);
  IV  NOT_10(G128,G712);
  IV  NOT_11(G139,G712);
  IV  NOT_12(G142,G29);
  IV  NOT_13(G143,G712);
  IV  NOT_14(G148,G712);
  IV  NOT_15(G153,G712);
  IV  NOT_16(G158,G712);
  IV  NOT_17(G165,G712);
  IV  NOT_18(G174,G712);
  IV  NOT_19(G176,G35);
  IV  NOT_20(G178,G34);
  IV  NOT_21(G179,G180);
  IV  NOT_22(G180,G92);
  IV  NOT_23(G188,G712);
  IV  NOT_24(G191,G36);
  IV  NOT_25(G192,G712);
  IV  NOT_26(G197,G712);
  IV  NOT_27(G204,G38);
  IV  NOT_28(G207,G712);
  IV  NOT_29(G210,G39);
  IV  NOT_30(G213,G712);
  IV  NOT_31(G216,G40);
  IV  NOT_32(G217,G712);
  IV  NOT_33(G236,G259);
  IV  NOT_34(G241,G259);
  IV  NOT_35(G246,G259);
  IV  NOT_36(G251,G259);
  IV  NOT_37(G258,G259);
  IV  NOT_38(G296,G297);
  IV  NOT_39(G302,G712);
  IV  NOT_40(G305,G324);
  IV  NOT_41(G308,G712);
  IV  NOT_42(G311,G324);
  IV  NOT_43(G314,G712);
  IV  NOT_44(G317,G324);
  IV  NOT_45(G320,G712);
  IV  NOT_46(G323,G324);
  IV  NOT_47(G336,G355);
  IV  NOT_48(G339,G355);
  IV  NOT_49(G343,G348);
  IV  NOT_50(G347,G348);
  IV  NOT_51(G348,G91);
  IV  NOT_52(G351,G645);
  IV  NOT_53(G354,G355);
  IV  NOT_54(G359,G372);
  IV  NOT_55(G364,G372);
  IV  NOT_56(G371,G372);
  IV  NOT_57(G378,G391);
  IV  NOT_58(G383,G391);
  IV  NOT_59(G390,G391);
  IV  NOT_60(G396,G404);
  IV  NOT_61(G403,G404);
  IV  NOT_62(G407,G712);
  IV  NOT_63(G415,G423);
  IV  NOT_64(G422,G423);
  IV  NOT_65(G426,G712);
  IV  NOT_66(G437,G712);
  IV  NOT_67(G440,G712);
  IV  NOT_68(G445,G65);
  IV  NOT_69(G446,G712);
  IV  NOT_70(G449,G66);
  IV  NOT_71(G450,G712);
  IV  NOT_72(G455,G456);
  IV  NOT_73(G458,G476);
  IV  NOT_74(G463,G476);
  IV  NOT_75(G468,G476);
  IV  NOT_76(G475,G476);
  IV  NOT_77(G486,G712);
  IV  NOT_78(G491,G500);
  IV  NOT_79(G495,G500);
  IV  NOT_80(G499,G500);
  IV  NOT_81(G504,G511);
  IV  NOT_82(G507,G511);
  IV  NOT_83(G510,G511);
  IV  NOT_84(G511,G63);
  IV  NOT_85(G525,G589);
  IV  NOT_86(G530,G589);
  IV  NOT_87(G535,G589);
  IV  NOT_88(G540,G589);
  IV  NOT_89(G547,G589);
  IV  NOT_90(G562,G610);
  IV  NOT_91(G566,G610);
  IV  NOT_92(G570,G610);
  IV  NOT_93(G574,G610);
  IV  NOT_94(G588,G589);
  IV  NOT_95(G595,G593);
  IV  NOT_96(G596,G597);
  IV  NOT_97(G600,G601);
  IV  NOT_98(G605,G610);
  IV  NOT_99(G609,G610);
  IV  NOT_100(G614,G64);
  IV  NOT_101(G615,G616);
  IV  NOT_102(G617,G645);
  IV  NOT_103(G620,G645);
  IV  NOT_104(G623,G645);
  IV  NOT_105(G626,G645);
  IV  NOT_106(G629,G645);
  IV  NOT_107(G632,G645);
  IV  NOT_108(G635,G645);
  IV  NOT_109(G638,G645);
  IV  NOT_110(G641,G645);
  IV  NOT_111(G644,G645);
  IV  NOT_112(G645,G90);
  IV  NOT_113(G656,G712);
  IV  NOT_114(G658,G659);
  IV  NOT_115(II1162,G13);
  IV  NOT_116(G659,II1162);
  IV  NOT_117(G661,G94);
  IV  NOT_118(G662,G712);
  IV  NOT_119(G665,G678);
  IV  NOT_120(G668,G712);
  IV  NOT_121(G671,G678);
  IV  NOT_122(G674,G712);
  IV  NOT_123(G677,G678);
  IV  NOT_124(II1183,G11);
  IV  NOT_125(G678,II1183);
  IV  NOT_126(G685,G696);
  IV  NOT_127(G689,G696);
  IV  NOT_128(G695,G696);
  IV  NOT_129(II1203,G10);
  IV  NOT_130(G696,II1203);
  IV  NOT_131(G701,G15);
  IV  NOT_132(II1211,G701);
  IV  NOT_133(G701BF,II1211);
  IV  NOT_134(G704,G712);
  IV  NOT_135(G706,G712);
  IV  NOT_136(G711,G712);
  IV  NOT_137(G712,G14);
  IV  NOT_138(G714,G701);
  IV  NOT_139(II1227,G6);
  IV  NOT_140(G715,II1227);
  IV  NOT_141(II1230,G7);
  IV  NOT_142(G716,II1230);
  IV  NOT_143(II1233,G8);
  IV  NOT_144(G717,II1233);
  IV  NOT_145(II1236,G9);
  IV  NOT_146(G718,II1236);
  IV  NOT_147(II1239,G12);
  IV  NOT_148(G719,II1239);
  IV  NOT_149(II1242,G0);
  IV  NOT_150(G720,II1242);
  IV  NOT_151(II1245,G1);
  IV  NOT_152(G721,II1245);
  IV  NOT_153(II1248,G2);
  IV  NOT_154(G722,II1248);
  IV  NOT_155(II1251,G3);
  IV  NOT_156(G723,II1251);
  IV  NOT_157(II1254,G4);
  IV  NOT_158(G724,II1254);
  IV  NOT_159(II1257,G5);
  IV  NOT_160(G725,II1257);
  IV  NOT_161(II1260,G93);
  IV  NOT_162(G726,II1260);
  IV  NOT_163(II1264,G16);
  IV  NOT_164(G728,II1264);
  IV  NOT_165(II1267,G95);
  IV  NOT_166(G729,II1267);
  AN2 AND2_0(G101,G630,G631);
  AN2 AND2_1(G102,G633,G634);
  AN2 AND2_2(G103,G636,G637);
  AN2 AND2_3(G104,G639,G640);
  AN2 AND2_4(G105,G642,G643);
  AN2 AND2_5(G109,G106,G108);
  AN2 AND2_6(G113,G114,G112);
  AN2 AND2_7(G116,G133,G25);
  AN2 AND2_8(G118,G119,G117);
  AN2 AND2_9(G121,G134,G26);
  AN2 AND2_10(G125,G122,G124);
  AN2 AND2_11(G129,G130,G128);
  AN2 AND2_12(G132,G136,G28);
  AN2 AND2_13(G133,G700,G111);
  AN2 AND2_14(G134,G133,G25);
  AN2 AND2_15(G135,G134,G26);
  AN2 AND2_16(G136,G135,G127);
  AN2 AND2_17(G140,G137,G139);
  AN2 AND2_18(G144,G145,G143);
  AN2 AND2_19(G147,G168,G30);
  AN2 AND2_20(G149,G150,G148);
  AN2 AND2_21(G152,G169,G31);
  AN2 AND2_22(G154,G155,G153);
  AN2 AND2_23(G157,G170,G32);
  AN2 AND2_24(G159,G160,G158);
  AN2 AND2_25(G162,G171,G33);
  AN2 AND2_26(G166,G163,G165);
  AN2 AND2_27(G168,G177,G142);
  AN2 AND2_28(G169,G168,G30);
  AN2 AND2_29(G170,G169,G31);
  AN2 AND2_30(G171,G170,G32);
  AN2 AND2_31(G172,G171,G33);
  AN2 AND2_32(G173,G172,G34);
  AN2 AND2_33(G175,G176,G174);
  AN2 AND2_34(G185,G181,G182);
  AN2 AND2_35(G189,G186,G188);
  AN2 AND2_36(G193,G194,G192);
  AN2 AND2_37(G196,G202,G37);
  AN2 AND2_38(G198,G199,G197);
  AN2 AND2_39(G201,G203,G38);
  AN2 AND2_40(G202,G522,G191);
  AN2 AND2_41(G203,G202,G37);
  AN2 AND2_42(G208,G205,G207);
  AN2 AND2_43(G214,G211,G213);
  AN2 AND2_44(G218,G219,G217);
  AN2 AND2_45(G221,G223,G41);
  AN2 AND2_46(G222,G183,G210);
  AN2 AND2_47(G223,G222,G216);
  AN2 AND2_48(G224,G203,G38);
  AN2 AND2_49(G225,G204,G203);
  AN2 AND2_50(G226,G136,G28);
  AN2 AND2_51(G227,G172,G178);
  AN2 AND2_52(G228,G223,G41);
  AN2 AND2_53(G229,G432,G62);
  AN2 AND2_54(G237,G238,G236);
  AN2 AND2_55(G240,G299,G42);
  AN2 AND2_56(G242,G243,G241);
  AN2 AND2_57(G245,G262,G43);
  AN2 AND2_58(G247,G248,G246);
  AN2 AND2_59(G250,G263,G44);
  AN2 AND2_60(G252,G253,G251);
  AN2 AND2_61(G255,G264,G45);
  AN2 AND2_62(G259,G624,G625);
  AN2 AND2_63(G260,G256,G258);
  AN2 AND2_64(G261,G265,G46);
  AN2 AND2_65(G262,G299,G42);
  AN2 AND2_66(G263,G262,G43);
  AN2 AND2_67(G264,G263,G44);
  AN2 AND2_68(G265,G264,G45);
  AN2 AND2_69(G271,G275,G266);
  AN2 AND2_70(G272,G276,G277);
  AN2 AND2_71(G273,G278,G279);
  AN2 AND2_72(G274,G280,G281);
  AN2 AND2_73(G303,G304,G302);
  AN2 AND2_74(G304,G306,G307);
  AN2 AND2_75(G309,G310,G308);
  AN2 AND2_76(G310,G312,G313);
  AN2 AND2_77(G315,G316,G314);
  AN2 AND2_78(G316,G318,G319);
  AN2 AND2_79(G321,G322,G320);
  AN2 AND2_80(G322,G325,G326);
  AN2 AND2_81(G329,G331,G714);
  AN2 AND2_82(G330,G332,G714);
  AN2 AND2_83(G335,G337,G338);
  AN2 AND2_84(G342,G344,G345);
  AN2 AND2_85(G346,G349,G350);
  AN2 AND2_86(G358,G523,G53);
  AN2 AND2_87(G360,G361,G359);
  AN2 AND2_88(G363,G523,G51);
  AN2 AND2_89(G365,G366,G364);
  AN2 AND2_90(G368,G375,G52);
  AN2 AND2_91(G373,G369,G371);
  AN2 AND2_92(G374,G376,G53);
  AN2 AND2_93(G375,G523,G51);
  AN2 AND2_94(G376,G375,G52);
  AN3 AND3_0(G377,G183,G54,G56);
  AN2 AND2_95(G379,G380,G378);
  AN2 AND2_96(G382,G183,G54);
  AN2 AND2_97(G384,G385,G383);
  AN2 AND2_98(G387,G394,G55);
  AN2 AND2_99(G392,G388,G390);
  AN2 AND2_100(G393,G395,G56);
  AN2 AND2_101(G394,G183,G54);
  AN2 AND2_102(G395,G394,G55);
  AN2 AND2_103(G397,G398,G396);
  AN2 AND2_104(G400,G335,G57);
  AN2 AND2_105(G405,G401,G403);
  AN2 AND2_106(G406,G412,G58);
  AN2 AND2_107(G408,G409,G407);
  AN2 AND2_108(G411,G413,G59);
  AN2 AND2_109(G412,G335,G57);
  AN2 AND2_110(G413,G335,G58);
  AN2 AND2_111(G414,G413,G59);
  AN2 AND2_112(G416,G417,G415);
  AN2 AND2_113(G419,G358,G60);
  AN2 AND2_114(G424,G420,G422);
  AN2 AND2_115(G425,G431,G61);
  AN2 AND2_116(G427,G428,G426);
  AN2 AND2_117(G430,G432,G62);
  AN2 AND2_118(G431,G358,G60);
  AN2 AND2_119(G432,G358,G61);
  AN2 AND2_120(G433,G356,G357);
  AN2 AND2_121(G435,G340,G341);
  AN2 AND2_122(G436,G352,G353);
  AN2 AND2_123(G438,G439,G437);
  AN2 AND2_124(G441,G442,G440);
  AN2 AND2_125(G443,G615,G511);
  AN2 AND2_126(G447,G448,G446);
  AN2 AND2_127(G451,G452,G450);
  AN2 AND2_128(G453,G615,G445);
  AN3 AND3_1(G457,G455,G449,G728);
  AN2 AND2_129(G459,G460,G458);
  AN2 AND2_130(G462,G434,G67);
  AN2 AND2_131(G464,G465,G463);
  AN2 AND2_132(G467,G479,G68);
  AN2 AND2_133(G469,G470,G468);
  AN2 AND2_134(G472,G480,G69);
  AN2 AND2_135(G477,G473,G475);
  AN2 AND2_136(G478,G481,G70);
  AN2 AND2_137(G479,G434,G67);
  AN2 AND2_138(G480,G479,G68);
  AN2 AND2_139(G481,G480,G69);
  AN2 AND2_140(G488,G505,G506);
  AN2 AND2_141(G489,G508,G509);
  AN2 AND2_142(G490,G512,G513);
  AN2 AND2_143(G494,G492,G493);
  AN2 AND2_144(G498,G496,G497);
  AN2 AND2_145(G503,G501,G502);
  AN2 AND2_146(G526,G527,G525);
  AN2 AND2_147(G529,G604,G74);
  AN2 AND2_148(G531,G532,G530);
  AN2 AND2_149(G534,G550,G75);
  AN2 AND2_150(G536,G537,G535);
  AN2 AND2_151(G539,G551,G76);
  AN2 AND2_152(G541,G542,G540);
  AN2 AND2_153(G544,G552,G77);
  AN2 AND2_154(G548,G545,G547);
  AN2 AND2_155(G549,G553,G78);
  AN2 AND2_156(G550,G604,G74);
  AN2 AND2_157(G551,G550,G75);
  AN2 AND2_158(G552,G551,G76);
  AN2 AND2_159(G553,G552,G77);
  AN2 AND2_160(G565,G563,G564);
  AN2 AND2_161(G569,G567,G568);
  AN2 AND2_162(G573,G571,G572);
  AN2 AND2_163(G577,G575,G576);
  AN2 AND2_164(G589,G627,G628);
  AN2 AND2_165(G590,G591,G588);
  AN2 AND2_166(G592,G594,G595);
  AN2 AND2_167(G601,G621,G622);
  AN2 AND2_168(G604,G433,G524);
  AN2 AND2_169(G608,G606,G607);
  AN2 AND2_170(G613,G611,G612);
  AN2 AND2_171(G648,G646,G647);
  AN2 AND2_172(G649,G618,G619);
  AN2 AND2_173(G650,G226,G661);
  AN2 AND2_174(G651,G227,G87);
  AN2 AND2_175(G652,G228,G88);
  AN2 AND2_176(G653,G229,G89);
  AN2 AND2_177(G654,G90,G476);
  AN2 AND2_178(G655,G91,G476);
  AN2 AND2_179(G657,G659,G656);
  AN2 AND2_180(G663,G664,G662);
  AN2 AND2_181(G664,G666,G667);
  AN2 AND2_182(G669,G670,G668);
  AN2 AND2_183(G670,G672,G673);
  AN2 AND2_184(G675,G676,G674);
  AN2 AND2_185(G676,G679,G680);
  AN2 AND2_186(G683,G684,G685);
  AN2 AND2_187(G688,G690,G691);
  AN2 AND2_188(G694,G697,G698);
  AN2 AND2_189(G702,G703,G645);
  AN2 AND2_190(G705,G230,G704);
  AN2 AND2_191(G707,G708,G706);
  AN2 AND2_192(G709,G678,G89);
  AN2 AND2_193(G713,G599,G711);
  AN2 AND2_194(G727,G476,G645);
  OR2 OR2_0(G110,G700,G111);
  OR2 OR2_1(G126,G135,G127);
  OR2 OR2_2(G141,G177,G142);
  OR2 OR2_3(G167,G172,G178);
  OR2 OR2_4(G177,G180,G226);
  OR2 OR2_5(G181,G178,G180);
  OR2 OR2_6(G182,G35,G179);
  OR2 OR2_7(G183,G180,G227);
  OR2 OR2_8(G184,G180,G173);
  OR2 OR2_9(G190,G522,G191);
  OR2 OR2_10(G209,G183,G210);
  OR2 OR2_11(G215,G222,G216);
  OR2 OR2_12(G235,G649,G233);
  OR2 OR2_13(G275,G101,G42);
  OR2 OR2_14(G276,G102,G43);
  OR2 OR2_15(G277,G267,G271);
  OR2 OR2_16(G278,G103,G44);
  OR2 OR2_17(G279,G268,G272);
  OR2 OR2_18(G280,G104,G45);
  OR2 OR2_19(G281,G269,G273);
  OR2 OR2_20(G282,G105,G46);
  OR2 OR2_21(G283,G270,G274);
  OR2 OR2_22(G291,G42,G101);
  OR2 OR2_23(G292,G43,G102);
  OR2 OR2_24(G293,G44,G103);
  OR2 OR2_25(G294,G45,G104);
  OR2 OR2_26(G295,G46,G105);
  OR4 OR4_0(G300,G50,G49,G48,G47);
  OR2 OR2_27(G306,G47,G324);
  OR2 OR2_28(G307,G719,G305);
  OR2 OR2_29(G312,G48,G324);
  OR2 OR2_30(G313,G47,G311);
  OR2 OR2_31(G318,G49,G324);
  OR2 OR2_32(G319,G48,G317);
  OR2 OR2_33(G324,G377,G348);
  OR2 OR2_34(G325,G50,G324);
  OR2 OR2_35(G326,G49,G323);
  OR2 OR2_36(G333,G300,G714);
  OR2 OR2_37(G334,G301,G714);
  OR2 OR2_38(G337,G224,G355);
  OR2 OR2_39(G338,G183,G336);
  OR2 OR2_40(G340,G38,G355);
  OR2 OR2_41(G341,G185,G339);
  OR2 OR2_42(G344,G229,G348);
  OR2 OR2_43(G345,G414,G343);
  OR2 OR2_44(G349,G62,G348);
  OR2 OR2_45(G350,G59,G347);
  OR2 OR2_46(G352,G346,G645);
  OR2 OR2_47(G353,G35,G351);
  OR2 OR2_48(G355,G457,G645);
  OR2 OR2_49(G356,G225,G355);
  OR2 OR2_50(G357,G184,G354);
  OR2 OR2_51(G372,G712,G358);
  OR2 OR2_52(G391,G712,G377);
  OR2 OR2_53(G404,G712,G413);
  OR2 OR2_54(G423,G712,G432);
  OR2 OR2_55(G434,G342,G645);
  OR2 OR2_56(G439,G435,G63);
  OR2 OR2_57(G448,G615,G65);
  OR2 OR2_58(G456,G83,G524);
  OR2 OR2_59(G492,G71,G500);
  OR2 OR2_60(G493,G488,G491);
  OR2 OR2_61(G496,G72,G500);
  OR2 OR2_62(G497,G489,G495);
  OR2 OR2_63(G500,G654,G712);
  OR2 OR2_64(G501,G73,G500);
  OR2 OR2_65(G502,G490,G499);
  OR2 OR2_66(G505,G723,G511);
  OR2 OR2_67(G506,G720,G504);
  OR2 OR2_68(G508,G724,G511);
  OR2 OR2_69(G509,G721,G507);
  OR2 OR2_70(G512,G725,G511);
  OR2 OR2_71(G513,G722,G510);
  OR2 OR2_72(G518,G71,G67);
  OR2 OR2_73(G519,G72,G68);
  OR2 OR2_74(G520,G73,G69);
  OR2 OR2_75(G521,G487,G70);
  OR2 OR2_76(G522,G348,G228);
  OR2 OR2_77(G523,G348,G414);
  OR2 OR2_78(G524,G554,G555);
  OR2 OR2_79(G563,G79,G610);
  OR2 OR2_80(G564,G715,G562);
  OR2 OR2_81(G567,G80,G610);
  OR2 OR2_82(G568,G716,G566);
  OR2 OR2_83(G571,G81,G610);
  OR2 OR2_84(G572,G717,G570);
  OR2 OR2_85(G575,G82,G610);
  OR2 OR2_86(G576,G718,G574);
  OR2 OR2_87(G583,G79,G74);
  OR2 OR2_88(G584,G80,G75);
  OR2 OR2_89(G585,G81,G76);
  OR2 OR2_90(G586,G82,G77);
  OR2 OR2_91(G587,G561,G78);
  OR2 OR2_92(G591,G592,G604);
  OR2 OR2_93(G594,G83,G593);
  OR2 OR2_94(G602,G85,G601);
  OR2 OR2_95(G603,G600,G84);
  OR2 OR2_96(G606,G84,G610);
  OR2 OR2_97(G607,G696,G605);
  OR2 OR2_98(G610,G655,G712);
  OR2 OR2_99(G611,G85,G610);
  OR2 OR2_100(G612,G678,G609);
  OR2 OR2_101(G618,G457,G645);
  OR2 OR2_102(G619,G715,G617);
  OR2 OR2_103(G621,G614,G645);
  OR2 OR2_104(G622,G717,G620);
  OR2 OR2_105(G624,G476,G645);
  OR2 OR2_106(G625,G716,G623);
  OR2 OR2_107(G627,G476,G645);
  OR2 OR2_108(G628,G718,G626);
  OR2 OR2_109(G630,G96,G645);
  OR2 OR2_110(G631,G720,G629);
  OR2 OR2_111(G633,G97,G645);
  OR2 OR2_112(G634,G721,G632);
  OR2 OR2_113(G636,G98,G645);
  OR2 OR2_114(G637,G722,G635);
  OR2 OR2_115(G639,G99,G645);
  OR2 OR2_116(G640,G723,G638);
  OR2 OR2_117(G642,G100,G645);
  OR2 OR2_118(G643,G724,G641);
  OR2 OR2_119(G646,G456,G645);
  OR2 OR2_120(G647,G725,G644);
  OR2 OR2_121(G666,G87,G678);
  OR2 OR2_122(G667,G661,G665);
  OR2 OR2_123(G672,G88,G678);
  OR2 OR2_124(G673,G87,G671);
  OR2 OR2_125(G679,G89,G678);
  OR2 OR2_126(G680,G88,G677);
  OR2 OR2_127(G682,G681,G699);
  OR2 OR2_128(G684,G645,G696);
  OR2 OR2_129(G687,G686,G699);
  OR2 OR2_130(G690,G348,G696);
  OR2 OR2_131(G691,G645,G689);
  OR2 OR2_132(G693,G692,G699);
  OR2 OR2_133(G697,G180,G696);
  OR2 OR2_134(G698,G348,G695);
  OR2 OR2_135(G699,G658,G712);
  ND2 NAND2_0(G96,G74,G596);
  ND2 NAND2_1(G97,G75,G596);
  ND2 NAND2_2(G98,G76,G596);
  ND2 NAND2_3(G99,G77,G596);
  ND2 NAND2_4(G100,G78,G596);
  ND2 NAND2_5(G106,G107,G110);
  ND2 NAND2_6(G107,G700,G111);
  ND2 NAND2_7(G122,G123,G126);
  ND2 NAND2_8(G123,G135,G127);
  ND2 NAND2_9(G137,G138,G141);
  ND2 NAND2_10(G138,G177,G142);
  ND2 NAND2_11(G163,G164,G167);
  ND2 NAND2_12(G164,G172,G178);
  ND2 NAND2_13(G186,G187,G190);
  ND2 NAND2_14(G187,G522,G191);
  ND2 NAND2_15(G205,G206,G209);
  ND2 NAND2_16(G206,G183,G210);
  ND2 NAND2_17(G211,G212,G215);
  ND2 NAND2_18(G212,G222,G216);
  ND2 NAND2_19(G230,G234,G235);
  ND2 NAND2_20(G231,G435,G648);
  ND3 NAND3_0(G232,G296,G298,G435);
  ND3 NAND3_1(G233,G700,G232,G231);
  ND2 NAND2_21(G234,G649,G436);
  ND2 NAND2_22(G266,G286,G291);
  ND2 NAND2_23(G267,G287,G292);
  ND2 NAND2_24(G268,G288,G293);
  ND2 NAND2_25(G269,G284,G294);
  ND2 NAND2_26(G270,G285,G295);
  ND2 NAND2_27(G284,G45,G104);
  ND2 NAND2_28(G285,G46,G105);
  ND2 NAND2_29(G286,G42,G101);
  ND2 NAND2_30(G287,G43,G102);
  ND2 NAND2_31(G288,G44,G103);
  ND2 NAND2_32(G297,G289,G290);
  ND2 NAND2_33(G298,G297,G700);
  ND4 NAND4_0(G301,G50,G49,G48,G47);
  ND2 NAND2_34(G331,G333,G22);
  ND2 NAND2_35(G332,G334,G331);
  ND2 NAND2_36(G476,G486,G616);
  ND2 NAND2_37(G482,G514,G518);
  ND2 NAND2_38(G483,G515,G519);
  ND2 NAND2_39(G484,G516,G520);
  ND2 NAND2_40(G485,G517,G521);
  ND2 NAND2_41(G514,G71,G67);
  ND2 NAND2_42(G515,G72,G68);
  ND2 NAND2_43(G516,G73,G69);
  ND2 NAND2_44(G517,G487,G70);
  ND3 NAND3_2(G554,G556,G557,G558);
  ND2 NAND2_45(G555,G559,G560);
  ND2 NAND2_46(G556,G578,G583);
  ND2 NAND2_47(G557,G579,G584);
  ND2 NAND2_48(G558,G580,G585);
  ND2 NAND2_49(G559,G581,G586);
  ND2 NAND2_50(G560,G582,G587);
  ND2 NAND2_51(G578,G79,G74);
  ND2 NAND2_52(G579,G80,G75);
  ND2 NAND2_53(G580,G81,G76);
  ND2 NAND2_54(G581,G82,G77);
  ND2 NAND2_55(G582,G561,G78);
  ND2 NAND2_56(G597,G602,G603);
  ND2 NAND2_57(G598,G435,G83);
  ND4 NAND4_1(G616,G482,G483,G484,G485);
  ND2 NAND2_58(G700,G282,G283);
  NR2 NOR2_0(G114,G115,G116);
  NR2 NOR2_1(G115,G133,G25);
  NR2 NOR2_2(G119,G120,G121);
  NR2 NOR2_3(G120,G134,G26);
  NR2 NOR2_4(G130,G131,G132);
  NR2 NOR2_5(G131,G136,G28);
  NR2 NOR2_6(G145,G146,G147);
  NR2 NOR2_7(G146,G168,G30);
  NR2 NOR2_8(G150,G151,G152);
  NR2 NOR2_9(G151,G169,G31);
  NR2 NOR2_10(G155,G156,G157);
  NR2 NOR2_11(G156,G170,G32);
  NR2 NOR2_12(G160,G161,G162);
  NR2 NOR2_13(G161,G171,G33);
  NR2 NOR2_14(G194,G195,G196);
  NR2 NOR2_15(G195,G202,G37);
  NR2 NOR2_16(G199,G200,G201);
  NR2 NOR2_17(G200,G203,G38);
  NR2 NOR2_18(G219,G220,G221);
  NR2 NOR2_19(G220,G223,G41);
  NR2 NOR2_20(G238,G239,G240);
  NR2 NOR2_21(G239,G299,G42);
  NR2 NOR2_22(G243,G244,G245);
  NR2 NOR2_23(G244,G262,G43);
  NR2 NOR2_24(G248,G249,G250);
  NR2 NOR2_25(G249,G263,G44);
  NR2 NOR2_26(G253,G254,G255);
  NR2 NOR2_27(G254,G264,G45);
  NR2 NOR2_28(G256,G257,G261);
  NR2 NOR2_29(G257,G265,G46);
  NR3 NOR3_0(G289,G270,G269,G268);
  NR2 NOR2_30(G290,G267,G266);
  NR2 NOR2_31(G299,G301,G328);
  NR2 NOR2_32(G327,G330,G23);
  NR2 NOR2_33(G328,G329,G327);
  NR2 NOR2_34(G361,G362,G363);
  NR2 NOR2_35(G362,G523,G51);
  NR2 NOR2_36(G366,G367,G368);
  NR2 NOR2_37(G367,G375,G52);
  NR2 NOR2_38(G369,G370,G374);
  NR2 NOR2_39(G370,G376,G53);
  NR2 NOR2_40(G380,G381,G382);
  NR2 NOR2_41(G381,G183,G54);
  NR2 NOR2_42(G385,G386,G387);
  NR2 NOR2_43(G386,G394,G55);
  NR2 NOR2_44(G388,G389,G393);
  NR2 NOR2_45(G389,G395,G56);
  NR2 NOR2_46(G398,G399,G400);
  NR2 NOR2_47(G399,G335,G57);
  NR2 NOR2_48(G401,G402,G406);
  NR2 NOR2_49(G402,G412,G58);
  NR2 NOR2_50(G409,G410,G411);
  NR2 NOR2_51(G410,G413,G59);
  NR2 NOR2_52(G417,G418,G419);
  NR2 NOR2_53(G418,G358,G60);
  NR2 NOR2_54(G420,G421,G425);
  NR2 NOR2_55(G421,G431,G61);
  NR2 NOR2_56(G428,G429,G430);
  NR2 NOR2_57(G429,G432,G62);
  NR2 NOR2_58(G442,G443,G444);
  NR2 NOR2_59(G444,G615,G64);
  NR2 NOR2_60(G452,G453,G454);
  NR2 NOR2_61(G454,G615,G66);
  NR2 NOR2_62(G460,G461,G462);
  NR2 NOR2_63(G461,G434,G67);
  NR2 NOR2_64(G465,G466,G467);
  NR2 NOR2_65(G466,G479,G68);
  NR2 NOR2_66(G470,G471,G472);
  NR2 NOR2_67(G471,G480,G69);
  NR2 NOR2_68(G473,G474,G478);
  NR2 NOR2_69(G474,G481,G70);
  NR3 NOR3_1(G487,G71,G72,G73);
  NR2 NOR2_70(G527,G528,G529);
  NR2 NOR2_71(G528,G604,G74);
  NR2 NOR2_72(G532,G533,G534);
  NR2 NOR2_73(G533,G550,G75);
  NR2 NOR2_74(G537,G538,G539);
  NR2 NOR2_75(G538,G551,G76);
  NR2 NOR2_76(G542,G543,G544);
  NR2 NOR2_77(G543,G552,G77);
  NR2 NOR2_78(G545,G546,G549);
  NR2 NOR2_79(G546,G553,G78);
  NR4 NOR4_0(G561,G79,G80,G81,G82);
  NR2 NOR2_80(G593,G435,G524);
  NR2 NOR2_81(G599,G598,G597);
  NR2 NOR2_82(G660,G658,G86);
  NR2 NOR2_83(G681,G683,G660);
  NR2 NOR2_84(G686,G688,G660);
  NR2 NOR2_85(G692,G694,G660);
  NR4 NOR4_1(G703,G650,G651,G652,G653);
  NR2 NOR2_86(G708,G709,G710);
  NR2 NOR2_87(G710,G678,G94);

endmodule
