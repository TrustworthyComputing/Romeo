module s5378(VDD,CK,n3065gat,n3066gat,n3067gat,n3068gat,n3069gat,n3070gat,
  n3071gat,
  n3072gat,n3073gat,n3074gat,n3075gat,n3076gat,n3077gat,n3078gat,n3079gat,
  n3080gat,n3081gat,n3082gat,n3083gat,n3084gat,n3085gat,n3086gat,n3087gat,
  n3088gat,n3089gat,n3090gat,n3091gat,n3092gat,n3093gat,n3094gat,n3095gat,
  n3097gat,n3098gat,n3099gat,n3100gat,n3104gat,n3105gat,n3106gat,n3107gat,
  n3108gat,n3109gat,n3110gat,n3111gat,n3112gat,n3113gat,n3114gat,n3115gat,
  n3116gat,n3117gat,n3118gat,n3119gat,n3120gat,n3121gat,n3122gat,n3123gat,
  n3124gat,n3125gat,n3126gat,n3127gat,n3128gat,n3129gat,n3130gat,n3131gat,
  n3132gat,n3133gat,n3134gat,n3135gat,n3136gat,n3137gat,n3138gat,n3139gat,
  n3140gat,n3141gat,n3142gat,n3143gat,n3144gat,n3145gat,n3146gat,n3147gat,
  n3148gat,n3149gat,n3150gat,n3151gat,n3152gat);
input VDD,CK,n3065gat,n3066gat,n3067gat,n3068gat,n3069gat,n3070gat,
  n3071gat,n3072gat,
  n3073gat,n3074gat,n3075gat,n3076gat,n3077gat,n3078gat,n3079gat,n3080gat,
  n3081gat,n3082gat,n3083gat,n3084gat,n3085gat,n3086gat,n3087gat,n3088gat,
  n3089gat,n3090gat,n3091gat,n3092gat,n3093gat,n3094gat,n3095gat,n3097gat,
  n3098gat,n3099gat,n3100gat;
output n3104gat,n3105gat,n3106gat,n3107gat,n3108gat,n3109gat,n3110gat,n3111gat,
  n3112gat,n3113gat,n3114gat,n3115gat,n3116gat,n3117gat,n3118gat,n3119gat,
  n3120gat,n3121gat,n3122gat,n3123gat,n3124gat,n3125gat,n3126gat,n3127gat,
  n3128gat,n3129gat,n3130gat,n3131gat,n3132gat,n3133gat,n3134gat,n3135gat,
  n3136gat,n3137gat,n3138gat,n3139gat,n3140gat,n3141gat,n3142gat,n3143gat,
  n3144gat,n3145gat,n3146gat,n3147gat,n3148gat,n3149gat,n3150gat,n3151gat,
  n3152gat;

  wire n673gat,n2897gat,n398gat,n2782gat,n402gat,n2790gat,n919gat,n2670gat,
    n846gat,n2793gat,n394gat,n703gat,n722gat,n726gat,n2510gat,n748gat,n271gat,
    n2732gat,n160gat,n2776gat,n337gat,n2735gat,n842gat,n2673gat,n341gat,
    n2779gat,n2522gat,n43gat,n2472gat,n1620gat,n2319gat,n2470gat,n1821gat,
    n1827gat,n1825gat,n2029gat,n1816gat,n1829gat,n2027gat,n283gat,n165gat,
    n279gat,n1026gat,n275gat,n2476gat,n55gat,n1068gat,n2914gat,n957gat,
    n2928gat,n861gat,n2927gat,n1294gat,n2896gat,n1241gat,n2922gat,n1298gat,
    n865gat,n2894gat,n1080gat,n2921gat,n1148gat,n2895gat,n2468gat,n933gat,
    n618gat,n491gat,n622gat,n626gat,n834gat,n3064gat,n707gat,n3055gat,n838gat,
    n3063gat,n830gat,n3062gat,n614gat,n3056gat,n2526gat,n504gat,n680gat,
    n2913gat,n816gat,n2920gat,n580gat,n2905gat,n824gat,n3057gat,n820gat,
    n3059gat,n883gat,n3058gat,n584gat,n2898gat,n684gat,n3060gat,n699gat,
    n3061gat,n2464gat,n567gat,n2399gat,n3048gat,n2343gat,n3049gat,n2203gat,
    n3051gat,n2562gat,n3047gat,n2207gat,n3050gat,n2626gat,n3040gat,n2490gat,
    n3044gat,n2622gat,n3042gat,n2630gat,n3037gat,n2543gat,n3041gat,n2102gat,
    n1606gat,n1880gat,n3052gat,n1763gat,n1610gat,n2155gat,n1858gat,n1035gat,
    n2918gat,n1121gat,n2952gat,n1072gat,n2919gat,n1282gat,n2910gat,n1226gat,
    n2907gat,n931gat,n2911gat,n1135gat,n2912gat,n1045gat,n2909gat,n1197gat,
    n2908gat,n2518gat,n2971gat,n667gat,n2904gat,n659gat,n2891gat,n553gat,
    n2903gat,n777gat,n2915gat,n561gat,n2901gat,n366gat,n2890gat,n322gat,
    n2888gat,n318gat,n2887gat,n314gat,n2886gat,n2599gat,n3010gat,n2588gat,
    n3016gat,n2640gat,n3054gat,n2658gat,n2579gat,n2495gat,n3036gat,n2390gat,
    n3034gat,n2270gat,n3031gat,n2339gat,n3035gat,n2502gat,n2646gat,n2634gat,
    n3053gat,n2506gat,n2613gat,n1834gat,n1625gat,n1767gat,n1626gat,n2084gat,
    n1603gat,n2143gat,n2541gat,n2061gat,n2557gat,n2139gat,n2487gat,n1899gat,
    n2532gat,n1850gat,n2628gat,n2403gat,n2397gat,n2394gat,n2341gat,n2440gat,
    n2560gat,n2407gat,n2205gat,n2347gat,n2201gat,n1389gat,n1793gat,n2021gat,
    n1781gat,n1394gat,n1516gat,n1496gat,n1392gat,n2091gat,n1685gat,n1332gat,
    n1565gat,n1740gat,n1330gat,n2179gat,n1945gat,n2190gat,n2268gat,n2135gat,
    n2337gat,n2262gat,n2388gat,n2182gat,n1836gat,n1433gat,n2983gat,n1316gat,
    n1431gat,n1363gat,n1314gat,n1312gat,n1361gat,n1775gat,n1696gat,n1871gat,
    n2009gat,n2592gat,n1773gat,n1508gat,n1636gat,n1678gat,n1712gat,n2309gat,
    n3000gat,n2450gat,n2307gat,n2446gat,n2661gat,n2095gat,n827gat,n2176gat,
    n2093gat,n2169gat,n2174gat,n2454gat,n2163gat,n2040gat,n1777gat,n2044gat,
    n2015gat,n2037gat,n2042gat,n2025gat,n2017gat,n2099gat,n2023gat,n2266gat,
    n2493gat,n2033gat,n2035gat,n2110gat,n2031gat,n2125gat,n2108gat,n2121gat,
    n2123gat,n2117gat,n2119gat,n1975gat,n2632gat,n2644gat,n2638gat,n156gat,
    n612gat,n152gat,n705gat,n331gat,n822gat,n388gat,n881gat,n463gat,n818gat,
    n327gat,n682gat,n384gat,n697gat,n256gat,n836gat,n470gat,n828gat,n148gat,
    n832gat,n2458gat,n2590gat,n2514gat,n2456gat,n1771gat,n1613gat,n1336gat,
    n1391gat,n1748gat,n1927gat,n1675gat,n1713gat,n1807gat,n1717gat,n1340gat,
    n1567gat,n1456gat,n1564gat,n1525gat,n1632gat,n1462gat,n1915gat,n1596gat,
    n1800gat,n1588gat,n1593gat,II1,n2717gat,n2715gat,II5,n2725gat,n2723gat,
    n296gat,n421gat,II11,n2768gat,II14,n2767gat,n373gat,II18,n2671gat,n2669gat,
    II23,n2845gat,n2844gat,II27,n2668gat,II30,n2667gat,n856gat,II44,n672gat,
    II47,n2783gat,II50,n396gat,II62,n2791gat,II65,II76,n401gat,n1645gat,
    n1499gat,II81,II92,n918gat,n1553gat,n1616gat,II97,n2794gat,II100,II111,
    n845gat,n1559gat,n1614gat,n1643gat,n1641gat,n1651gat,n1642gat,n1562gat,
    n1556gat,n1560gat,n1557gat,n1640gat,n1639gat,n1566gat,n1605gat,n1554gat,
    n1555gat,n1722gat,n1558gat,n392gat,II149,n702gat,n1319gat,n1256gat,n720gat,
    II171,n725gat,n1447gat,n1117gat,n1627gat,n1618gat,II178,n721gat,n1380gat,
    n1114gat,n1628gat,n1621gat,n701gat,n1446gat,n1318gat,n1705gat,n1619gat,
    n1706gat,n1622gat,II192,n2856gat,n2854gat,II196,n1218gat,II199,n2861gat,
    n2859gat,II203,n1219gat,II206,n2864gat,n2862gat,II210,n1220gat,II214,
    n2860gat,II217,n1221gat,II220,n2863gat,II223,n1222gat,II227,n2855gat,II230,
    n1223gat,n640gat,n1213gat,II237,n753gat,II240,n2716gat,II243,n2869gat,
    n2867gat,II248,n2868gat,II253,n2906gat,n754gat,II256,n2724gat,II259,
    n2728gat,n2726gat,II264,n2727gat,n422gat,n2889gat,II270,n755gat,n747gat,
    II275,n756gat,II278,n757gat,II282,n758gat,n2508gat,II297,n2733gat,II300,
    II311,n270gat,II314,n263gat,II317,n2777gat,II320,II331,n159gat,II334,
    n264gat,II337,n2736gat,II340,II351,n336gat,II354,n265gat,n158gat,II359,
    n266gat,n335gat,II363,n267gat,n269gat,II368,n268gat,n41gat,n258gat,II375,
    n48gat,II378,n1018gat,II381,n2674gat,II384,II395,n841gat,II398,n1019gat,
    II401,n1020gat,n840gat,II406,n1021gat,II409,n1022gat,n724gat,II414,
    n1023gat,II420,n1013gat,n49gat,II423,n2780gat,II426,II437,n340gat,II440,
    n480gat,II443,n481gat,II446,n393gat,II449,n482gat,II453,n483gat,II456,
    n484gat,n339gat,II461,n485gat,n42gat,n475gat,II468,n50gat,n162gat,II473,
    n51gat,II476,n52gat,II480,n53gat,n2520gat,n1448gat,n1376gat,n1701gat,
    n1617gat,n1379gat,n1377gat,n1615gat,n1624gat,n1500gat,n1113gat,n1503gat,
    n1501gat,n1779gat,n1623gat,II509,n2730gat,II512,n2729gat,n2317gat,n1819gat,
    n1823gat,n1817gat,II572,n1828gat,II576,n2851gat,II579,n2850gat,II583,
    n2786gat,n2785gat,n92gat,n637gat,n529gat,n293gat,n361gat,II591,n2722gat,
    II594,n2721gat,n297gat,II606,n282gat,II609,n172gat,II620,n164gat,II623,
    n173gat,II634,n278gat,II637,n174gat,n163gat,II642,n175gat,n277gat,II646,
    n176gat,n281gat,II651,n177gat,n54gat,n167gat,II658,n60gat,II661,n911gat,
    II672,n1025gat,II675,n912gat,II678,n913gat,n1024gat,II683,n914gat,n917gat,
    II687,n915gat,n844gat,II692,n916gat,II698,n906gat,n61gat,II709,n274gat,
    II712,n348gat,II715,n349gat,II718,n397gat,II721,n350gat,n400gat,II726,
    n351gat,II729,n352gat,n273gat,II734,n353gat,n178gat,n343gat,II741,n62gat,
    n66gat,II746,n63gat,II749,n64gat,II753,n65gat,n2474gat,II768,n2832gat,
    II771,n2831gat,n2731gat,II776,n2719gat,n2718gat,II790,n1067gat,II793,
    n949gat,II796,n2839gat,n2838gat,n2775gat,II812,n956gat,II815,n950gat,II818,
    n2712gat,n2711gat,n2734gat,II834,n860gat,II837,n951gat,n955gat,II842,
    n952gat,n859gat,II846,n953gat,n1066gat,II851,n954gat,n857gat,n944gat,II858,
    n938gat,n2792gat,II863,n2847gat,n2846gat,II877,n1293gat,II880,n1233gat,
    n2672gat,II885,n2853gat,n2852gat,II899,n1240gat,II902,n1234gat,II913,
    n1297gat,II916,n1235gat,n1239gat,II921,n1236gat,n1296gat,II925,n1237gat,
    n1292gat,II930,n1238gat,II936,n1228gat,n939gat,n2778gat,II941,n2837gat,
    n2836gat,II955,n864gat,II958,n1055gat,n2789gat,II963,n2841gat,n2840gat,
    II977,n1079gat,II980,n1056gat,n2781gat,II985,n2843gat,n2842gat,II999,
    n1147gat,II1002,n1057gat,n1078gat,II1007,n1058gat,n1146gat,II1011,n1059gat,
    n863gat,II1016,n1060gat,n928gat,n1050gat,II1023,n940gat,n858gat,II1028,
    n941gat,II1031,n942gat,II1035,n943gat,n2466gat,n2720gat,n740gat,n2784gat,
    n743gat,n746gat,n294gat,n360gat,n374gat,n616gat,II1067,n501gat,n489gat,
    II1079,n502gat,II1082,n617gat,II1085,n499gat,II1088,n490gat,II1091,n500gat,
    n620gat,II1103,n738gat,n624gat,II1115,n737gat,II1118,n621gat,II1121,
    n733gat,II1124,n625gat,II1127,n735gat,II1138,n833gat,II1141,n714gat,II1152,
    n706gat,II1155,n715gat,II1166,n837gat,II1169,n716gat,II1174,n717gat,II1178,
    n718gat,II1183,n719gat,n515gat,n709gat,II1190,n509gat,II1201,n829gat,
    II1204,n734gat,II1209,n736gat,II1216,n728gat,n510gat,II1227,n613gat,II1230,
    n498gat,II1236,n503gat,n404gat,n493gat,II1243,n511gat,n405gat,II1248,
    n512gat,II1251,n513gat,II1255,n514gat,n2524gat,n17gat,n564gat,n79gat,
    n86gat,n219gat,n78gat,n563gat,II1278,n289gat,n179gat,n287gat,n188gat,
    n288gat,n72gat,n181gat,n111gat,n182gat,II1302,n679gat,II1305,n808gat,
    II1319,n815gat,II1322,n809gat,II1336,n579gat,II1339,n810gat,n814gat,II1344,
    n811gat,n578gat,II1348,n812gat,n678gat,II1353,n813gat,n677gat,n803gat,
    II1360,n572gat,II1371,n823gat,II1374,n591gat,II1385,n819gat,II1388,n592gat,
    II1399,n882gat,II1402,n593gat,II1407,n594gat,II1411,n595gat,II1416,n596gat,
    II1422,n586gat,n573gat,II1436,n583gat,II1439,n691gat,II1450,n683gat,II1453,
    n692gat,II1464,n698gat,II1467,n693gat,II1472,n694gat,II1476,n695gat,
    n582gat,II1481,n696gat,n456gat,n686gat,II1488,n574gat,n565gat,II1493,
    n575gat,II1496,n576gat,II1500,n577gat,n2462gat,n2665gat,II1516,n2596gat,
    n189gat,n286gat,n194gat,n187gat,n21gat,n15gat,II1538,n2398gat,n2353gat,
    II1550,n2342gat,n2284gat,n2354gat,n2356gat,n2214gat,n2286gat,II1585,
    n2624gat,II1606,n2489gat,II1617,n2621gat,n2533gat,n2534gat,II1630,n2629gat,
    n2486gat,n2429gat,n2432gat,n2430gat,II1655,n2101gat,n1693gat,II1667,
    n1879gat,n1698gat,n1934gat,n1543gat,II1683,n1762gat,n1673gat,n2989gat,
    II1698,n2154gat,n2488gat,II1703,n2625gat,n2530gat,n2531gat,II1708,n2542gat,
    n2482gat,n2426gat,n2480gat,n2153gat,n2355gat,II1719,n2561gat,n2443gat,
    n2289gat,II1724,n2148gat,II1734,n855gat,n759gat,II1749,n1034gat,II1752,
    n1189gat,n1075gat,II1766,n1120gat,II1769,n1190gat,n760gat,II1783,n1071gat,
    II1786,n1191gat,n1119gat,II1791,n1192gat,n1070gat,II1795,n1193gat,n1033gat,
    II1800,n1194gat,n1183gat,n1184gat,II1807,n1274gat,n644gat,n1280gat,n641gat,
    II1833,n1225gat,II1837,n1281gat,n1224gat,II1843,n2970gat,n1275gat,n761gat,
    II1857,n930gat,II1860,n1206gat,n762gat,II1874,n1134gat,II1877,n1207gat,
    n643gat,II1891,n1044gat,II1894,n1208gat,n1133gat,II1899,n1209gat,n1043gat,
    II1903,n1210gat,n929gat,II1908,n1211gat,n1268gat,n1201gat,II1915,n1276gat,
    n1329gat,II1920,n1277gat,II1923,n1278gat,II1927,n1279gat,n1284gat,n1269gat,
    n642gat,n1195gat,II1947,n1196gat,n2516gat,II1961,n3017gat,n851gat,n853gat,
    n1725gat,n664gat,n852gat,n854gat,II1981,n666gat,n368gat,II1996,n658gat,
    II1999,n784gat,n662gat,II2014,n552gat,II2017,n785gat,n661gat,II2032,
    n776gat,II2035,n786gat,n551gat,II2040,n787gat,n775gat,II2044,n788gat,
    n657gat,II2049,n789gat,n35gat,n779gat,II2056,n125gat,n558gat,n559gat,
    n371gat,II2084,n365gat,II2088,n560gat,n364gat,II2094,n2876gat,n126gat,
    n663gat,II2109,n321gat,II2112,n226gat,n370gat,II2127,n317gat,II2130,
    n227gat,n369gat,II2145,n313gat,II2148,n228gat,n316gat,II2153,n229gat,
    n312gat,II2157,n230gat,n320gat,II2162,n231gat,n34gat,n221gat,II2169,
    n127gat,n133gat,II2174,n128gat,II2177,n129gat,II2181,n130gat,n665gat,
    n1601gat,n120gat,n2597gat,n2595gat,n2594gat,n2586gat,II2213,n2573gat,
    II2225,n2574gat,II2228,n2575gat,II2232,n2639gat,II2235,n2576gat,II2238,
    n2577gat,II2242,n2578gat,II2248,n2568gat,n2582gat,II2251,n2206gat,II2254,
    n2414gat,II2257,n2415gat,II2260,n2202gat,II2263,n2416gat,II2268,n2417gat,
    II2271,n2418gat,II2275,n2419gat,II2281,n2409gat,n2585gat,n2656gat,II2316,
    n2389gat,II2319,n2494gat,II2324,n3014gat,n2649gat,II2344,n2338gat,II2349,
    n2269gat,II2354,n2880gat,n2652gat,n2500gat,n2620gat,n2612gat,II2372,
    n2606gat,II2376,n2607gat,n2540gat,II2380,n2608gat,n2536gat,II2385,n2609gat,
    II2389,n2610gat,II2394,n2611gat,II2400,n2601gat,n2616gat,II2403,n2550gat,
    II2414,n2633gat,II2417,n2551gat,II2420,n2552gat,II2425,n2553gat,II2428,
    n2554gat,II2433,n2555gat,II2439,n2545gat,n2619gat,n2504gat,n2660gat,
    n2655gat,n1528gat,n2293gat,n1523gat,n2219gat,n1592gat,n1529gat,n2666gat,
    n1704gat,n2422gat,n3013gat,n2290gat,n2081gat,n2218gat,n2285gat,n2359gat,
    n2358gat,n1414gat,n1415gat,n566gat,n1480gat,n2292gat,n1301gat,n1416gat,
    n1150gat,n873gat,n2011gat,n2306gat,n1478gat,n1481gat,n875gat,n1410gat,
    n2357gat,n876gat,n1347gat,n1160gat,n1484gat,n1084gat,n983gat,n1482gat,
    n2363gat,n1157gat,n1483gat,n985gat,n1530gat,n2364gat,n1307gat,n1308gat,
    n1085gat,n1479gat,n2291gat,n1348gat,n1349gat,n2217gat,n1591gat,n2223gat,
    n1437gat,n1438gat,n1832gat,n1765gat,n1878gat,n1442gat,n1831gat,n1444gat,
    n1378gat,n2975gat,n1322gat,n2974gat,n1439gat,n1486gat,n1370gat,n1426gat,
    n1369gat,n2966gat,n1366gat,n1365gat,n1374gat,n2979gat,n2162gat,n2220gat,
    n1450gat,n1423gat,n1427gat,n1608gat,n2082gat,n1449gat,n1494gat,n1590gat,
    n1248gat,n2954gat,n1418gat,n1417gat,n1306gat,n2964gat,n1353gat,n1419gat,
    n1247gat,n2958gat,n1355gat,n1422gat,n1300gat,n2963gat,n1487gat,n1485gat,
    n1164gat,n2953gat,n1356gat,n1354gat,n1436gat,n1435gat,n1106gat,n2949gat,
    n1425gat,n1421gat,n1105gat,n2934gat,n1424gat,n1420gat,n1309gat,n2959gat,
    II2672,n2142gat,n1788gat,II2684,n2060gat,n1786gat,II2696,n2138gat,n1839gat,
    n1897gat,n1884gat,n1848gat,n1783gat,n1548gat,II2721,n1719gat,n2137gat,
    n1633gat,n2059gat,n1785gat,II2731,n1849gat,n1784gat,n1716gat,II2736,
    n1635gat,n2401gat,n1989gat,n2392gat,n1918gat,II2771,n2439gat,n1986gat,
    n1866gat,n1865gat,II2785,n2406gat,n2216gat,n2345gat,n1988gat,n1735gat,
    n1861gat,n1387gat,n1694gat,II2813,n1780gat,n2019gat,n1549gat,II2832,
    n1551gat,II2837,n2346gat,n2152gat,n2405gat,n2351gat,II2843,n2402gat,
    n2212gat,II2847,n2393gat,n1991gat,n1665gat,n1666gat,n1517gat,n1578gat,
    II2873,n1495gat,n1604gat,II2885,n2090gat,n1550gat,II2890,n1552gat,n1738gat,
    II2915,n1739gat,n1925gat,n1920gat,n1917gat,n1921gat,n2141gat,n1787gat,
    II2926,n1859gat,n1922gat,n1798gat,II2935,n1743gat,n1923gat,n1864gat,
    n1690gat,II2953,n2178gat,n1661gat,n1660gat,n1572gat,n1576gat,n2438gat,
    n2283gat,n1520gat,n1582gat,n1580gat,n1577gat,n1990gat,n2988gat,II2978,
    n2189gat,II2989,n2134gat,II3000,n2261gat,n2128gat,n2129gat,n1695gat,II3016,
    n2181gat,II3056,n1311gat,n1707gat,n1659gat,n2987gat,n1515gat,n1521gat,
    n1736gat,n1737gat,n1658gat,n1724gat,n1732gat,n1662gat,n1663gat,n1656gat,
    n1655gat,n1670gat,n1667gat,n1569gat,n1570gat,n1568gat,n1575gat,n1727gat,
    n1728gat,n1797gat,n1801gat,n1730gat,n1731gat,n1561gat,n1571gat,n1668gat,
    n1734gat,n1742gat,n1671gat,n1669gat,n1652gat,n1657gat,n1648gat,n1729gat,
    n1790gat,n1726gat,n2004gat,n1929gat,n1869gat,II3143,n2591gat,n1584gat,
    n1714gat,II3149,n1718gat,II3163,n1507gat,n1396gat,n1401gat,II3168,n1393gat,
    n1409gat,n1476gat,II3174,n1898gat,n1838gat,II3179,II3191,n1677gat,n2000gat,
    n1412gat,n2001gat,n1999gat,II3211,n2663gat,n3018gat,n2448gat,n2662gat,
    n2444gat,II3235,n2238gat,n3019gat,n1310gat,n199gat,n87gat,n195gat,n184gat,
    n204gat,II3273,n2168gat,n2452gat,n1691gat,II3287,n3020gat,II3290,n3021gat,
    II3293,n3022gat,n1699gat,II3297,n3023gat,II3300,n3024gat,II3303,n3025gat,
    II3306,n3026gat,II3309,n3027gat,II3312,n3028gat,II3315,n3029gat,II3318,
    n3030gat,n2260gat,n2257gat,n2188gat,n2187gat,n3004gat,II3336,n2039gat,
    II3339,n1774gat,II3342,n1315gat,n2097gat,n1855gat,n2014gat,II3387,n2194gat,
    II3390,n3032gat,n2256gat,II3394,n3033gat,n2251gat,n2184gat,n3003gat,II3401,
    n2192gat,n2133gat,n2131gat,n2185gat,n2049gat,n3001gat,II3412,n2057gat,
    n2253gat,n2252gat,n2248gat,n3006gat,n2264gat,II3429,n2265gat,n2492gat,
    n2329gat,II3436,n1709gat,n1845gat,n1891gat,n1963gat,n1886gat,n1968gat,
    n1958gat,n1629gat,n1895gat,n1631gat,n1711gat,n2990gat,n2200gat,n2078gat,
    n2437gat,n2195gat,II3457,n2556gat,n1956gat,II3461,n3038gat,n1954gat,II3465,
    n3039gat,n1888gat,n2048gat,n2994gat,II3472,n2539gat,n1969gat,n1893gat,
    n1892gat,n2993gat,II3483,n2436gat,n2056gat,n2998gat,II3491,n2387gat,II3494,
    n3043gat,n1960gat,n1887gat,n1961gat,n2996gat,II3504,n2330gat,n2199gat,
    n2147gat,II3509,n3045gat,n2332gat,II3513,n3046gat,n2259gat,n2328gat,
    n3008gat,II3520,n2498gat,n2151gat,n2193gat,n2209gat,n3005gat,II3530,
    n2396gat,n2052gat,n2058gat,n2997gat,II3539,n2198gat,n2349gat,n2215gat,
    n2281gat,n3009gat,II3549,n2197gat,n2146gat,n3002gat,II3558,n2196gat,II3587,
    n2124gat,n2115gat,II3610,n1882gat,II3621,n1974gat,n1955gat,n1970gat,
    n1896gat,n1973gat,n2558gat,n2559gat,II3635,II3646,n2643gat,n2333gat,
    n2564gat,n2352gat,n2642gat,n2636gat,n2637gat,II3660,n88gat,n84gat,n375gat,
    n110gat,II3677,n155gat,n253gat,n1702gat,n150gat,II3691,n151gat,n243gat,
    n233gat,n154gat,n800gat,n2874gat,II3703,n2917gat,n235gat,n2878gat,II3713,
    n2892gat,n372gat,n212gat,n329gat,II3736,n387gat,n334gat,n1700gat,n386gat,
    II3742,n330gat,n1430gat,n1490gat,n452gat,n2885gat,II3754,n2900gat,n333gat,
    n2883gat,II3765,n2929gat,II3777,n462gat,n325gat,n457gat,n2884gat,n461gat,
    n458gat,n2902gat,II3801,n2925gat,n144gat,n247gat,II3808,n326gat,n878gat,
    n2879gat,II3817,n2916gat,n382gat,II3831,n383gat,n134gat,n2875gat,II3841,
    n2899gat,n254gat,n252gat,n2877gat,n468gat,II3867,n469gat,n381gat,n2893gat,
    II3876,n2926gat,n241gat,n140gat,II3882,n255gat,n802gat,n2882gat,II3891,
    n2924gat,n146gat,II3904,n147gat,n380gat,n2881gat,II3914,n2923gat,n69gat,
    n68gat,n1885gat,II3923,n2710gat,n2707gat,n16gat,n295gat,n357gat,n11gat,
    n12gat,n1889gat,II3935,n2704gat,n2700gat,n2051gat,II3941,n2684gat,n2680gat,
    n1350gat,II3945,n2696gat,II3948,n2692gat,II3951,n2683gat,II3954,n2679gat,
    II3957,n2449gat,n1754gat,II3962,n2830gat,n2827gat,n2512gat,n1544gat,
    n1769gat,n1683gat,n1756gat,n2167gat,n2013gat,II4000,n1791gat,n2691gat,
    n2695gat,n1518gat,n2699gat,n2703gat,n2159gat,n2478gat,II4014,n2744gat,
    n2740gat,n2158gat,n2186gat,II4020,n2800gat,n2797gat,n2288gat,II4024,
    n1513gat,n2537gat,n2538gat,n2442gat,n2483gat,n1334gat,II4055,n1747gat,
    II4067,n1674gat,n1403gat,n1402gat,II4081,n1806gat,n1634gat,n1338gat,II4105,
    n1455gat,II4108,n1339gat,n1505gat,n2980gat,II4117,n2758gat,n2755gat,
    n1546gat,II4122,n2752gat,n2748gat,n2012gat,n2016gat,n2002gat,n2008gat,
    II4129,n2858gat,n2857gat,II4135,n2766gat,II4138,n2765gat,n1684gat,n1759gat,
    II4145,II4157,n1524gat,n1862gat,n1863gat,n1919gat,n1860gat,n1460gat,II4185,
    n1595gat,n1454gat,n1469gat,n1468gat,n1519gat,II4194,n1461gat,n1477gat,
    n2984gat,n1594gat,II4212,n1587gat,n1681gat,II4217,II4222,n1761gat,n2751gat,
    n2747gat,II4227,n1760gat,n2743gat,n2739gat,n1978gat,II4233,n1721gat,
    n2808gat,II4236,n2804gat,n517gat,n518gat,n417gat,n418gat,n413gat,n411gat,
    n412gat,n522gat,n406gat,n516gat,n407gat,n355gat,n290gat,n525gat,n527gat,
    n356gat,n416gat,n415gat,n528gat,n521gat,n358gat,n532gat,n639gat,n523gat,
    n1111gat,n635gat,n524gat,n414gat,n1112gat,n630gat,n741gat,n629gat,n633gat,
    n634gat,n926gat,n632gat,n670gat,n636gat,n1123gat,n1007gat,n1006gat,II4309,
    n2941gat,n2814gat,II4312,n2811gat,n1002gat,n2946gat,II4329,n2950gat,
    n2813gat,II4332,n2810gat,n888gat,n2933gat,II4349,n2935gat,n2818gat,II4352,
    n2816gat,n898gat,n2940gat,II4369,n2937gat,n2817gat,II4372,n2815gat,
    n1179gat,n2947gat,II4389,n2956gat,n2824gat,II4392,n2821gat,n897gat,
    n2939gat,II4409,n2938gat,n2823gat,II4412,n2820gat,n894gat,n2932gat,II4429,
    n2936gat,n2829gat,II4432,n2826gat,n1180gat,n2948gat,II4449,n2955gat,
    n2828gat,II4452,n2825gat,n671gat,n628gat,n631gat,n976gat,II4475,n2951gat,
    n2807gat,II4478,n2803gat,n2127gat,II4482,n2682gat,II4485,n2678gat,n2046gat,
    II4489,n2681gat,II4492,n2677gat,n1708gat,II4496,n2688gat,II4499,n2686gat,
    n455gat,n291gat,n2237gat,II4506,n2764gat,n2763gat,n1782gat,II4512,n2762gat,
    n2760gat,n2325gat,II4518,n2761gat,n2759gat,n2245gat,II4524,n2757gat,
    n2754gat,n2244gat,II4530,n2756gat,n2753gat,n2243gat,II4536,n2750gat,
    n2746gat,n2246gat,II4542,n2749gat,n2745gat,n2384gat,II4548,n2742gat,
    n2738gat,n2385gat,II4554,n2741gat,n2737gat,n1286gat,II4558,n2687gat,
    n2685gat,n1328gat,n1381gat,n1384gat,II4566,n2694gat,n2690gat,n1382gat,
    n1451gat,n1453gat,II4573,n2693gat,n2689gat,n927gat,n925gat,n1452gat,II4580,
    n2702gat,n2698gat,n923gat,n921gat,n1890gat,II4587,n2701gat,n2697gat,
    n850gat,n739gat,n1841gat,II4594,n2709gat,n2706gat,n922gat,n848gat,n2047gat,
    II4601,n2708gat,n2705gat,n924gat,n849gat,n2050gat,II4608,n2799gat,n2796gat,
    n1118gat,n1032gat,n2054gat,II4615,n2798gat,n2795gat,II4620,n1745gat,
    n2806gat,II4623,n2802gat,II4626,n1870gat,n1086gat,II4630,n2805gat,II4633,
    n2801gat,n67gat,n85gat,n71gat,n180gat,n1840gat,II4642,n2812gat,n2809gat,
    n76gat,n82gat,n14gat,n186gat,n1842gat,II4651,n2822gat,n2819gat,II4654,
    II4657,II4660,II4663,II4666,II4669,II4672,II4675,II4678,II4681,II4684,
    II4687,II4690,II4693,II4696,II4699,II4702,II4705,II4708,II4711,II4714,
    II4717,II4720,II4723,II4726,II4729,II4732,II4735,II4738,II4741,II4744,
    II4747,II4750,II4753,II4756,II4759,II4762,II4765,II4768,II4771,II4774,
    II4777,II4780,II4783,II4786,II4789,II4792,II4795,II4798,n648gat,n442gat,
    n1214gat,n1215gat,n1216gat,n1217gat,n745gat,n638gat,n423gat,n362gat,
    n749gat,n750gat,n751gat,n752gat,n259gat,n260gat,n261gat,n262gat,n1014gat,
    n1015gat,n1016gat,n1017gat,n476gat,n477gat,n478gat,n479gat,n44gat,n45gat,
    n46gat,n47gat,n168gat,n169gat,n170gat,n171gat,n907gat,n908gat,n909gat,
    n910gat,n344gat,n345gat,n346gat,n347gat,n56gat,n57gat,n58gat,n59gat,
    n768gat,n655gat,n963gat,n868gat,n962gat,n959gat,n945gat,n946gat,n947gat,
    n948gat,n647gat,n441gat,n967gat,n792gat,n1229gat,n1230gat,n1231gat,
    n1232gat,n443gat,n439gat,n966gat,n790gat,n444gat,n440gat,n1051gat,n1052gat,
    n1053gat,n1054gat,n934gat,n935gat,n936gat,n937gat,n710gat,n711gat,n712gat,
    n713gat,n729gat,n730gat,n731gat,n732gat,n494gat,n495gat,n496gat,n497gat,
    n505gat,n506gat,n507gat,n508gat,II1277,n767gat,n653gat,n867gat,n771gat,
    n964gat,n961gat,n804gat,n805gat,n806gat,n807gat,n587gat,n588gat,n589gat,
    n590gat,n447gat,n445gat,n687gat,n688gat,n689gat,n690gat,n568gat,n569gat,
    n570gat,n571gat,II1515,II1584,n1692gat,II1723,II1733,n2428gat,n769gat,
    n1076gat,n766gat,n1185gat,n1186gat,n1187gat,n1188gat,n645gat,n646gat,
    n1383gat,n1327gat,n651gat,n652gat,n765gat,n1202gat,n1203gat,n1204gat,
    n1205gat,n1270gat,n1271gat,n1272gat,n1273gat,n763gat,n1287gat,n1285gat,
    n793gat,n556gat,n795gat,n656gat,n794gat,n773gat,n965gat,n960gat,n780gat,
    n781gat,n782gat,n783gat,n555gat,n450gat,n654gat,n557gat,n874gat,n132gat,
    n649gat,n449gat,n791gat,n650gat,n774gat,n764gat,n222gat,n223gat,n224gat,
    n225gat,n121gat,n122gat,n123gat,n124gat,n2460gat,n2423gat,n2569gat,
    n2570gat,n2571gat,n2572gat,n2410gat,n2411gat,n2412gat,n2413gat,n2580gat,
    n2581gat,n2567gat,n2499gat,n299gat,n207gat,n2647gat,n2648gat,n2602gat,
    n2603gat,n2604gat,n2605gat,n2546gat,n2547gat,n2548gat,n2549gat,n2614gat,
    n2615gat,n2461gat,n2421gat,n2930gat,n1153gat,n1151gat,n982gat,n877gat,
    n2957gat,n1159gat,n1158gat,n1156gat,n1155gat,n1443gat,n1325gat,n1321gat,
    n1320gat,n1368gat,n1258gat,n1373gat,n1372gat,n2978gat,n1441gat,n1440gat,
    n1371gat,n1367gat,n2982gat,n1504gat,n1502gat,n1250gat,n1103gat,n1304gat,
    n1249gat,n1246gat,n1161gat,n1291gat,n1245gat,n2973gat,n1352gat,n1351gat,
    n1303gat,n1302gat,n1163gat,n1102gat,n1101gat,n996gat,n1104gat,n887gat,
    n1305gat,n1162gat,n2977gat,n1360gat,n1359gat,n1358gat,n1357gat,II2720,
    II2735,II2812,n1703gat,n1778gat,n1609gat,II2831,II2889,II2925,II2934,
    n1733gat,n1581gat,n2079gat,n2073gat,n1574gat,n1573gat,n2992gat,n1723gat,
    n1647gat,n1646gat,n2986gat,n1650gat,n1649gat,n1563gat,n2991gat,n1654gat,
    n1653gat,n1644gat,II3148,II3178,n2981gat,n1413gat,n1408gat,n1407gat,
    n2258gat,n2255gat,n2132gat,n2130gat,n3007gat,n2250gat,n2249gat,n1710gat,
    n1630gat,n1894gat,n1847gat,n1846gat,n2055gat,n1967gat,n1959gat,n1957gat,
    n2211gat,n2210gat,n2053gat,n1964gat,n2350gat,n2282gat,n2213gat,n2150gat,
    n2149gat,n2995gat,n1962gat,n2999gat,n1972gat,n1971gat,n3011gat,n2331gat,
    n3015gat,n2566gat,n2565gat,n141gat,n38gat,n37gat,n1074gat,n872gat,n234gat,
    n137gat,n378gat,n377gat,n250gat,n249gat,n248gat,n869gat,n453gat,n448gat,
    n251gat,n244gat,n974gat,n973gat,n870gat,n246gat,n245gat,n460gat,n459gat,
    n975gat,n972gat,n969gat,n145gat,n143gat,n971gat,n970gat,n968gat,n142gat,
    n40gat,n39gat,n772gat,n451gat,n446gat,n139gat,n136gat,n391gat,n390gat,
    n1083gat,n1077gat,n242gat,n240gat,n871gat,n797gat,n324gat,n238gat,n237gat,
    n1082gat,n796gat,n1599gat,II3999,n1586gat,n1755gat,II4023,n1470gat,
    n1400gat,n1399gat,n1398gat,II4144,n1467gat,n1466gat,n2985gat,n1686gat,
    n1533gat,n1532gat,n1531gat,II4216,n2931gat,n1100gat,n994gat,n989gat,
    n880gat,n2943gat,n1012gat,n905gat,n1003gat,n902gat,n1099gat,n998gat,
    n995gat,n980gat,n2960gat,n1175gat,n1174gat,n1001gat,n999gat,n2969gat,
    n1323gat,n1264gat,n981gat,n890gat,n889gat,n886gat,n892gat,n891gat,n2942gat,
    n904gat,n903gat,n1152gat,n1092gat,n997gat,n993gat,n900gat,n895gat,n1094gat,
    n1093gat,n988gat,n984gat,n2965gat,n1267gat,n1257gat,n1178gat,n1116gat,
    n2961gat,n1375gat,n1324gat,n1091gat,n1088gat,n992gat,n987gat,n899gat,
    n896gat,n2967gat,n1262gat,n1260gat,n1098gat,n1090gat,n986gat,n885gat,
    n901gat,n893gat,n1097gat,n1089gat,n1087gat,n991gat,n2968gat,n1326gat,
    n1261gat,n1177gat,n1115gat,n2944gat,n977gat,n2945gat,n1096gat,n1095gat,
    n990gat,n979gat,n2962gat,n1176gat,n1173gat,n1004gat,n1000gat,n1029gat,
    n1028gat,n1031gat,n1030gat,n1011gat,n1181gat,n1010gat,n1005gat,n1182gat,
    n73gat,n70gat,n77gat,n13gat,n1935gat,n197gat,n22gat,n93gat,n2239gat,
    n2433gat,n2427gat,n2583gat,n2650gat,n2617gat,n1598gat,n1154gat,n1411gat,
    n1498gat,n1607gat,n1428gat,n1794gat,n1796gat,n1792gat,n1406gat,n2664gat,
    n1926gat,n1916gat,n1994gat,n1924gat,n1758gat,n200gat,n196gat,n2018gat,
    n89gat,n1471gat,n1472gat,n1600gat,n1397gat,n2005gat,n1818gat,n1510gat,
    n1459gat,n1458gat,n1602gat,n520gat,n519gat,n410gat,n354gat,n408gat,n526gat,
    n531gat,n530gat,n359gat,n420gat,n801gat,n879gat,n1255gat,n1009gat,n409gat,
    n292gat,n419gat,n1243gat,n1171gat,n1244gat,n1265gat,n1254gat,n1008gat,
    n1253gat,n1266gat,n1200gat,n1172gat,n1251gat,n1259gat,n1212gat,n1263gat,
    n978gat,n1199gat,n1252gat,n1757gat;

  FD1 DFF_0(CK,n673gat,n2897gat);
  FD1 DFF_1(CK,n398gat,n2782gat);
  FD1 DFF_2(CK,n402gat,n2790gat);
  FD1 DFF_3(CK,n919gat,n2670gat);
  FD1 DFF_4(CK,n846gat,n2793gat);
  FD1 DFF_5(CK,n394gat,n2782gat);
  FD1 DFF_6(CK,n703gat,n2790gat);
  FD1 DFF_7(CK,n722gat,n2670gat);
  FD1 DFF_8(CK,n726gat,n2793gat);
  FD1 DFF_9(CK,n2510gat,n748gat);
  FD1 DFF_10(CK,n271gat,n2732gat);
  FD1 DFF_11(CK,n160gat,n2776gat);
  FD1 DFF_12(CK,n337gat,n2735gat);
  FD1 DFF_13(CK,n842gat,n2673gat);
  FD1 DFF_14(CK,n341gat,n2779gat);
  FD1 DFF_15(CK,n2522gat,n43gat);
  FD1 DFF_16(CK,n2472gat,n1620gat);
  FD1 DFF_17(CK,n2319gat,n2470gat);
  FD1 DFF_18(CK,n1821gat,n1827gat);
  FD1 DFF_19(CK,n1825gat,n1827gat);
  FD1 DFF_20(CK,n2029gat,n1816gat);
  FD1 DFF_21(CK,n1829gat,n2027gat);
  FD1 DFF_22(CK,n283gat,n2732gat);
  FD1 DFF_23(CK,n165gat,n2776gat);
  FD1 DFF_24(CK,n279gat,n2735gat);
  FD1 DFF_25(CK,n1026gat,n2673gat);
  FD1 DFF_26(CK,n275gat,n2779gat);
  FD1 DFF_27(CK,n2476gat,n55gat);
  FD1 DFF_28(CK,n1068gat,n2914gat);
  FD1 DFF_29(CK,n957gat,n2928gat);
  FD1 DFF_30(CK,n861gat,n2927gat);
  FD1 DFF_31(CK,n1294gat,n2896gat);
  FD1 DFF_32(CK,n1241gat,n2922gat);
  FD1 DFF_33(CK,n1298gat,n2897gat);
  FD1 DFF_34(CK,n865gat,n2894gat);
  FD1 DFF_35(CK,n1080gat,n2921gat);
  FD1 DFF_36(CK,n1148gat,n2895gat);
  FD1 DFF_37(CK,n2468gat,n933gat);
  FD1 DFF_38(CK,n618gat,n2790gat);
  FD1 DFF_39(CK,n491gat,n2782gat);
  FD1 DFF_40(CK,n622gat,n2793gat);
  FD1 DFF_41(CK,n626gat,n2670gat);
  FD1 DFF_42(CK,n834gat,n3064gat);
  FD1 DFF_43(CK,n707gat,n3055gat);
  FD1 DFF_44(CK,n838gat,n3063gat);
  FD1 DFF_45(CK,n830gat,n3062gat);
  FD1 DFF_46(CK,n614gat,n3056gat);
  FD1 DFF_47(CK,n2526gat,n504gat);
  FD1 DFF_48(CK,n680gat,n2913gat);
  FD1 DFF_49(CK,n816gat,n2920gat);
  FD1 DFF_50(CK,n580gat,n2905gat);
  FD1 DFF_51(CK,n824gat,n3057gat);
  FD1 DFF_52(CK,n820gat,n3059gat);
  FD1 DFF_53(CK,n883gat,n3058gat);
  FD1 DFF_54(CK,n584gat,n2898gat);
  FD1 DFF_55(CK,n684gat,n3060gat);
  FD1 DFF_56(CK,n699gat,n3061gat);
  FD1 DFF_57(CK,n2464gat,n567gat);
  FD1 DFF_58(CK,n2399gat,n3048gat);
  FD1 DFF_59(CK,n2343gat,n3049gat);
  FD1 DFF_60(CK,n2203gat,n3051gat);
  FD1 DFF_61(CK,n2562gat,n3047gat);
  FD1 DFF_62(CK,n2207gat,n3050gat);
  FD1 DFF_63(CK,n2626gat,n3040gat);
  FD1 DFF_64(CK,n2490gat,n3044gat);
  FD1 DFF_65(CK,n2622gat,n3042gat);
  FD1 DFF_66(CK,n2630gat,n3037gat);
  FD1 DFF_67(CK,n2543gat,n3041gat);
  FD1 DFF_68(CK,n2102gat,n1606gat);
  FD1 DFF_69(CK,n1880gat,n3052gat);
  FD1 DFF_70(CK,n1763gat,n1610gat);
  FD1 DFF_71(CK,n2155gat,n1858gat);
  FD1 DFF_72(CK,n1035gat,n2918gat);
  FD1 DFF_73(CK,n1121gat,n2952gat);
  FD1 DFF_74(CK,n1072gat,n2919gat);
  FD1 DFF_75(CK,n1282gat,n2910gat);
  FD1 DFF_76(CK,n1226gat,n2907gat);
  FD1 DFF_77(CK,n931gat,n2911gat);
  FD1 DFF_78(CK,n1135gat,n2912gat);
  FD1 DFF_79(CK,n1045gat,n2909gat);
  FD1 DFF_80(CK,n1197gat,n2908gat);
  FD1 DFF_81(CK,n2518gat,n2971gat);
  FD1 DFF_82(CK,n667gat,n2904gat);
  FD1 DFF_83(CK,n659gat,n2891gat);
  FD1 DFF_84(CK,n553gat,n2903gat);
  FD1 DFF_85(CK,n777gat,n2915gat);
  FD1 DFF_86(CK,n561gat,n2901gat);
  FD1 DFF_87(CK,n366gat,n2890gat);
  FD1 DFF_88(CK,n322gat,n2888gat);
  FD1 DFF_89(CK,n318gat,n2887gat);
  FD1 DFF_90(CK,n314gat,n2886gat);
  FD1 DFF_91(CK,n2599gat,n3010gat);
  FD1 DFF_92(CK,n2588gat,n3016gat);
  FD1 DFF_93(CK,n2640gat,n3054gat);
  FD1 DFF_94(CK,n2658gat,n2579gat);
  FD1 DFF_95(CK,n2495gat,n3036gat);
  FD1 DFF_96(CK,n2390gat,n3034gat);
  FD1 DFF_97(CK,n2270gat,n3031gat);
  FD1 DFF_98(CK,n2339gat,n3035gat);
  FD1 DFF_99(CK,n2502gat,n2646gat);
  FD1 DFF_100(CK,n2634gat,n3053gat);
  FD1 DFF_101(CK,n2506gat,n2613gat);
  FD1 DFF_102(CK,n1834gat,n1625gat);
  FD1 DFF_103(CK,n1767gat,n1626gat);
  FD1 DFF_104(CK,n2084gat,n1603gat);
  FD1 DFF_105(CK,n2143gat,n2541gat);
  FD1 DFF_106(CK,n2061gat,n2557gat);
  FD1 DFF_107(CK,n2139gat,n2487gat);
  FD1 DFF_108(CK,n1899gat,n2532gat);
  FD1 DFF_109(CK,n1850gat,n2628gat);
  FD1 DFF_110(CK,n2403gat,n2397gat);
  FD1 DFF_111(CK,n2394gat,n2341gat);
  FD1 DFF_112(CK,n2440gat,n2560gat);
  FD1 DFF_113(CK,n2407gat,n2205gat);
  FD1 DFF_114(CK,n2347gat,n2201gat);
  FD1 DFF_115(CK,n1389gat,n1793gat);
  FD1 DFF_116(CK,n2021gat,n1781gat);
  FD1 DFF_117(CK,n1394gat,n1516gat);
  FD1 DFF_118(CK,n1496gat,n1392gat);
  FD1 DFF_119(CK,n2091gat,n1685gat);
  FD1 DFF_120(CK,n1332gat,n1565gat);
  FD1 DFF_121(CK,n1740gat,n1330gat);
  FD1 DFF_122(CK,n2179gat,n1945gat);
  FD1 DFF_123(CK,n2190gat,n2268gat);
  FD1 DFF_124(CK,n2135gat,n2337gat);
  FD1 DFF_125(CK,n2262gat,n2388gat);
  FD1 DFF_126(CK,n2182gat,n1836gat);
  FD1 DFF_127(CK,n1433gat,n2983gat);
  FD1 DFF_128(CK,n1316gat,n1431gat);
  FD1 DFF_129(CK,n1363gat,n1314gat);
  FD1 DFF_130(CK,n1312gat,n1361gat);
  FD1 DFF_131(CK,n1775gat,n1696gat);
  FD1 DFF_132(CK,n1871gat,n2009gat);
  FD1 DFF_133(CK,n2592gat,n1773gat);
  FD1 DFF_134(CK,n1508gat,n1636gat);
  FD1 DFF_135(CK,n1678gat,n1712gat);
  FD1 DFF_136(CK,n2309gat,n3000gat);
  FD1 DFF_137(CK,n2450gat,n2307gat);
  FD1 DFF_138(CK,n2446gat,n2661gat);
  FD1 DFF_139(CK,n2095gat,n827gat);
  FD1 DFF_140(CK,n2176gat,n2093gat);
  FD1 DFF_141(CK,n2169gat,n2174gat);
  FD1 DFF_142(CK,n2454gat,n2163gat);
  FD1 DFF_143(CK,n2040gat,n1777gat);
  FD1 DFF_144(CK,n2044gat,n2015gat);
  FD1 DFF_145(CK,n2037gat,n2042gat);
  FD1 DFF_146(CK,n2025gat,n2017gat);
  FD1 DFF_147(CK,n2099gat,n2023gat);
  FD1 DFF_148(CK,n2266gat,n2493gat);
  FD1 DFF_149(CK,n2033gat,n2035gat);
  FD1 DFF_150(CK,n2110gat,n2031gat);
  FD1 DFF_151(CK,n2125gat,n2108gat);
  FD1 DFF_152(CK,n2121gat,n2123gat);
  FD1 DFF_153(CK,n2117gat,n2119gat);
  FD1 DFF_154(CK,n1975gat,n2632gat);
  FD1 DFF_155(CK,n2644gat,n2638gat);
  FD1 DFF_156(CK,n156gat,n612gat);
  FD1 DFF_157(CK,n152gat,n705gat);
  FD1 DFF_158(CK,n331gat,n822gat);
  FD1 DFF_159(CK,n388gat,n881gat);
  FD1 DFF_160(CK,n463gat,n818gat);
  FD1 DFF_161(CK,n327gat,n682gat);
  FD1 DFF_162(CK,n384gat,n697gat);
  FD1 DFF_163(CK,n256gat,n836gat);
  FD1 DFF_164(CK,n470gat,n828gat);
  FD1 DFF_165(CK,n148gat,n832gat);
  FD1 DFF_166(CK,n2458gat,n2590gat);
  FD1 DFF_167(CK,n2514gat,n2456gat);
  FD1 DFF_168(CK,n1771gat,n1613gat);
  FD1 DFF_169(CK,n1336gat,n1391gat);
  FD1 DFF_170(CK,n1748gat,n1927gat);
  FD1 DFF_171(CK,n1675gat,n1713gat);
  FD1 DFF_172(CK,n1807gat,n1717gat);
  FD1 DFF_173(CK,n1340gat,n1567gat);
  FD1 DFF_174(CK,n1456gat,n1564gat);
  FD1 DFF_175(CK,n1525gat,n1632gat);
  FD1 DFF_176(CK,n1462gat,n1915gat);
  FD1 DFF_177(CK,n1596gat,n1800gat);
  FD1 DFF_178(CK,n1588gat,n1593gat);
  IV  NOT_0(II1,n3088gat);
  IV  NOT_1(n2717gat,II1);
  IV  NOT_2(n2715gat,n2717gat);
  IV  NOT_3(II5,n3087gat);
  IV  NOT_4(n2725gat,II5);
  IV  NOT_5(n2723gat,n2725gat);
  IV  NOT_6(n296gat,n421gat);
  IV  NOT_7(II11,n3093gat);
  IV  NOT_8(n2768gat,II11);
  IV  NOT_9(II14,n2768gat);
  IV  NOT_10(n2767gat,II14);
  IV  NOT_11(n373gat,n2767gat);
  IV  NOT_12(II18,n3072gat);
  IV  NOT_13(n2671gat,II18);
  IV  NOT_14(n2669gat,n2671gat);
  IV  NOT_15(II23,n3081gat);
  IV  NOT_16(n2845gat,II23);
  IV  NOT_17(n2844gat,n2845gat);
  IV  NOT_18(II27,n3095gat);
  IV  NOT_19(n2668gat,II27);
  IV  NOT_20(II30,n2668gat);
  IV  NOT_21(n2667gat,II30);
  IV  NOT_22(n856gat,n2667gat);
  IV  NOT_23(II44,n673gat);
  IV  NOT_24(n672gat,II44);
  IV  NOT_25(II47,n3069gat);
  IV  NOT_26(n2783gat,II47);
  IV  NOT_27(II50,n2783gat);
  IV  NOT_28(n2782gat,II50);
  IV  NOT_29(n396gat,n398gat);
  IV  NOT_30(II62,n3070gat);
  IV  NOT_31(n2791gat,II62);
  IV  NOT_32(II65,n2791gat);
  IV  NOT_33(n2790gat,II65);
  IV  NOT_34(II76,n402gat);
  IV  NOT_35(n401gat,II76);
  IV  NOT_36(n1645gat,n1499gat);
  IV  NOT_37(II81,n2671gat);
  IV  NOT_38(n2670gat,II81);
  IV  NOT_39(II92,n919gat);
  IV  NOT_40(n918gat,II92);
  IV  NOT_41(n1553gat,n1616gat);
  IV  NOT_42(II97,n3071gat);
  IV  NOT_43(n2794gat,II97);
  IV  NOT_44(II100,n2794gat);
  IV  NOT_45(n2793gat,II100);
  IV  NOT_46(II111,n846gat);
  IV  NOT_47(n845gat,II111);
  IV  NOT_48(n1559gat,n1614gat);
  IV  NOT_49(n1643gat,n1641gat);
  IV  NOT_50(n1651gat,n1642gat);
  IV  NOT_51(n1562gat,n1556gat);
  IV  NOT_52(n1560gat,n1557gat);
  IV  NOT_53(n1640gat,n1639gat);
  IV  NOT_54(n1566gat,n1605gat);
  IV  NOT_55(n1554gat,n1555gat);
  IV  NOT_56(n1722gat,n1558gat);
  IV  NOT_57(n392gat,n394gat);
  IV  NOT_58(II149,n703gat);
  IV  NOT_59(n702gat,II149);
  IV  NOT_60(n1319gat,n1256gat);
  IV  NOT_61(n720gat,n722gat);
  IV  NOT_62(II171,n726gat);
  IV  NOT_63(n725gat,II171);
  IV  NOT_64(n1447gat,n1117gat);
  IV  NOT_65(n1627gat,n1618gat);
  IV  NOT_66(II178,n722gat);
  IV  NOT_67(n721gat,II178);
  IV  NOT_68(n1380gat,n1114gat);
  IV  NOT_69(n1628gat,n1621gat);
  IV  NOT_70(n701gat,n703gat);
  IV  NOT_71(n1446gat,n1318gat);
  IV  NOT_72(n1705gat,n1619gat);
  IV  NOT_73(n1706gat,n1622gat);
  IV  NOT_74(II192,n3083gat);
  IV  NOT_75(n2856gat,II192);
  IV  NOT_76(n2854gat,n2856gat);
  IV  NOT_77(II196,n2854gat);
  IV  NOT_78(n1218gat,II196);
  IV  NOT_79(II199,n3085gat);
  IV  NOT_80(n2861gat,II199);
  IV  NOT_81(n2859gat,n2861gat);
  IV  NOT_82(II203,n2859gat);
  IV  NOT_83(n1219gat,II203);
  IV  NOT_84(II206,n3084gat);
  IV  NOT_85(n2864gat,II206);
  IV  NOT_86(n2862gat,n2864gat);
  IV  NOT_87(II210,n2862gat);
  IV  NOT_88(n1220gat,II210);
  IV  NOT_89(II214,n2861gat);
  IV  NOT_90(n2860gat,II214);
  IV  NOT_91(II217,n2860gat);
  IV  NOT_92(n1221gat,II217);
  IV  NOT_93(II220,n2864gat);
  IV  NOT_94(n2863gat,II220);
  IV  NOT_95(II223,n2863gat);
  IV  NOT_96(n1222gat,II223);
  IV  NOT_97(II227,n2856gat);
  IV  NOT_98(n2855gat,II227);
  IV  NOT_99(II230,n2855gat);
  IV  NOT_100(n1223gat,II230);
  IV  NOT_101(n640gat,n1213gat);
  IV  NOT_102(II237,n640gat);
  IV  NOT_103(n753gat,II237);
  IV  NOT_104(II240,n2717gat);
  IV  NOT_105(n2716gat,II240);
  IV  NOT_106(II243,n3089gat);
  IV  NOT_107(n2869gat,II243);
  IV  NOT_108(n2867gat,n2869gat);
  IV  NOT_109(II248,n2869gat);
  IV  NOT_110(n2868gat,II248);
  IV  NOT_111(II253,n2906gat);
  IV  NOT_112(n754gat,II253);
  IV  NOT_113(II256,n2725gat);
  IV  NOT_114(n2724gat,II256);
  IV  NOT_115(II259,n3086gat);
  IV  NOT_116(n2728gat,II259);
  IV  NOT_117(n2726gat,n2728gat);
  IV  NOT_118(II264,n2728gat);
  IV  NOT_119(n2727gat,II264);
  IV  NOT_120(n422gat,n2889gat);
  IV  NOT_121(II270,n422gat);
  IV  NOT_122(n755gat,II270);
  IV  NOT_123(n747gat,n2906gat);
  IV  NOT_124(II275,n747gat);
  IV  NOT_125(n756gat,II275);
  IV  NOT_126(II278,n2889gat);
  IV  NOT_127(n757gat,II278);
  IV  NOT_128(II282,n1213gat);
  IV  NOT_129(n758gat,II282);
  IV  NOT_130(n2508gat,n2510gat);
  IV  NOT_131(II297,n3065gat);
  IV  NOT_132(n2733gat,II297);
  IV  NOT_133(II300,n2733gat);
  IV  NOT_134(n2732gat,II300);
  IV  NOT_135(II311,n271gat);
  IV  NOT_136(n270gat,II311);
  IV  NOT_137(II314,n270gat);
  IV  NOT_138(n263gat,II314);
  IV  NOT_139(II317,n3067gat);
  IV  NOT_140(n2777gat,II317);
  IV  NOT_141(II320,n2777gat);
  IV  NOT_142(n2776gat,II320);
  IV  NOT_143(II331,n160gat);
  IV  NOT_144(n159gat,II331);
  IV  NOT_145(II334,n159gat);
  IV  NOT_146(n264gat,II334);
  IV  NOT_147(II337,n3066gat);
  IV  NOT_148(n2736gat,II337);
  IV  NOT_149(II340,n2736gat);
  IV  NOT_150(n2735gat,II340);
  IV  NOT_151(II351,n337gat);
  IV  NOT_152(n336gat,II351);
  IV  NOT_153(II354,n336gat);
  IV  NOT_154(n265gat,II354);
  IV  NOT_155(n158gat,n160gat);
  IV  NOT_156(II359,n158gat);
  IV  NOT_157(n266gat,II359);
  IV  NOT_158(n335gat,n337gat);
  IV  NOT_159(II363,n335gat);
  IV  NOT_160(n267gat,II363);
  IV  NOT_161(n269gat,n271gat);
  IV  NOT_162(II368,n269gat);
  IV  NOT_163(n268gat,II368);
  IV  NOT_164(n41gat,n258gat);
  IV  NOT_165(II375,n41gat);
  IV  NOT_166(n48gat,II375);
  IV  NOT_167(II378,n725gat);
  IV  NOT_168(n1018gat,II378);
  IV  NOT_169(II381,n3073gat);
  IV  NOT_170(n2674gat,II381);
  IV  NOT_171(II384,n2674gat);
  IV  NOT_172(n2673gat,II384);
  IV  NOT_173(II395,n842gat);
  IV  NOT_174(n841gat,II395);
  IV  NOT_175(II398,n841gat);
  IV  NOT_176(n1019gat,II398);
  IV  NOT_177(II401,n721gat);
  IV  NOT_178(n1020gat,II401);
  IV  NOT_179(n840gat,n842gat);
  IV  NOT_180(II406,n840gat);
  IV  NOT_181(n1021gat,II406);
  IV  NOT_182(II409,n720gat);
  IV  NOT_183(n1022gat,II409);
  IV  NOT_184(n724gat,n726gat);
  IV  NOT_185(II414,n724gat);
  IV  NOT_186(n1023gat,II414);
  IV  NOT_187(II420,n1013gat);
  IV  NOT_188(n49gat,II420);
  IV  NOT_189(II423,n3068gat);
  IV  NOT_190(n2780gat,II423);
  IV  NOT_191(II426,n2780gat);
  IV  NOT_192(n2779gat,II426);
  IV  NOT_193(II437,n341gat);
  IV  NOT_194(n340gat,II437);
  IV  NOT_195(II440,n340gat);
  IV  NOT_196(n480gat,II440);
  IV  NOT_197(II443,n702gat);
  IV  NOT_198(n481gat,II443);
  IV  NOT_199(II446,n394gat);
  IV  NOT_200(n393gat,II446);
  IV  NOT_201(II449,n393gat);
  IV  NOT_202(n482gat,II449);
  IV  NOT_203(II453,n701gat);
  IV  NOT_204(n483gat,II453);
  IV  NOT_205(II456,n392gat);
  IV  NOT_206(n484gat,II456);
  IV  NOT_207(n339gat,n341gat);
  IV  NOT_208(II461,n339gat);
  IV  NOT_209(n485gat,II461);
  IV  NOT_210(n42gat,n475gat);
  IV  NOT_211(II468,n42gat);
  IV  NOT_212(n50gat,II468);
  IV  NOT_213(n162gat,n1013gat);
  IV  NOT_214(II473,n162gat);
  IV  NOT_215(n51gat,II473);
  IV  NOT_216(II476,n475gat);
  IV  NOT_217(n52gat,II476);
  IV  NOT_218(II480,n258gat);
  IV  NOT_219(n53gat,II480);
  IV  NOT_220(n2520gat,n2522gat);
  IV  NOT_221(n1448gat,n1376gat);
  IV  NOT_222(n1701gat,n1617gat);
  IV  NOT_223(n1379gat,n1377gat);
  IV  NOT_224(n1615gat,n1624gat);
  IV  NOT_225(n1500gat,n1113gat);
  IV  NOT_226(n1503gat,n1501gat);
  IV  NOT_227(n1779gat,n1623gat);
  IV  NOT_228(II509,n3099gat);
  IV  NOT_229(n2730gat,II509);
  IV  NOT_230(II512,n2730gat);
  IV  NOT_231(n2729gat,II512);
  IV  NOT_232(n2470gat,n2472gat);
  IV  NOT_233(n2317gat,n2319gat);
  IV  NOT_234(n1819gat,n1821gat);
  IV  NOT_235(n1823gat,n1825gat);
  IV  NOT_236(n1816gat,n1817gat);
  IV  NOT_237(n2027gat,n2029gat);
  IV  NOT_238(II572,n1829gat);
  IV  NOT_239(n1828gat,II572);
  IV  NOT_240(II576,n3100gat);
  IV  NOT_241(n2851gat,II576);
  IV  NOT_242(II579,n2851gat);
  IV  NOT_243(n2850gat,II579);
  IV  NOT_244(II583,n2786gat);
  IV  NOT_245(n2785gat,II583);
  IV  NOT_246(n92gat,n2785gat);
  IV  NOT_247(n637gat,n529gat);
  IV  NOT_248(n293gat,n361gat);
  IV  NOT_249(II591,n3094gat);
  IV  NOT_250(n2722gat,II591);
  IV  NOT_251(II594,n2722gat);
  IV  NOT_252(n2721gat,II594);
  IV  NOT_253(n297gat,n2721gat);
  IV  NOT_254(II606,n283gat);
  IV  NOT_255(n282gat,II606);
  IV  NOT_256(II609,n282gat);
  IV  NOT_257(n172gat,II609);
  IV  NOT_258(II620,n165gat);
  IV  NOT_259(n164gat,II620);
  IV  NOT_260(II623,n164gat);
  IV  NOT_261(n173gat,II623);
  IV  NOT_262(II634,n279gat);
  IV  NOT_263(n278gat,II634);
  IV  NOT_264(II637,n278gat);
  IV  NOT_265(n174gat,II637);
  IV  NOT_266(n163gat,n165gat);
  IV  NOT_267(II642,n163gat);
  IV  NOT_268(n175gat,II642);
  IV  NOT_269(n277gat,n279gat);
  IV  NOT_270(II646,n277gat);
  IV  NOT_271(n176gat,II646);
  IV  NOT_272(n281gat,n283gat);
  IV  NOT_273(II651,n281gat);
  IV  NOT_274(n177gat,II651);
  IV  NOT_275(n54gat,n167gat);
  IV  NOT_276(II658,n54gat);
  IV  NOT_277(n60gat,II658);
  IV  NOT_278(II661,n845gat);
  IV  NOT_279(n911gat,II661);
  IV  NOT_280(II672,n1026gat);
  IV  NOT_281(n1025gat,II672);
  IV  NOT_282(II675,n1025gat);
  IV  NOT_283(n912gat,II675);
  IV  NOT_284(II678,n918gat);
  IV  NOT_285(n913gat,II678);
  IV  NOT_286(n1024gat,n1026gat);
  IV  NOT_287(II683,n1024gat);
  IV  NOT_288(n914gat,II683);
  IV  NOT_289(n917gat,n919gat);
  IV  NOT_290(II687,n917gat);
  IV  NOT_291(n915gat,II687);
  IV  NOT_292(n844gat,n846gat);
  IV  NOT_293(II692,n844gat);
  IV  NOT_294(n916gat,II692);
  IV  NOT_295(II698,n906gat);
  IV  NOT_296(n61gat,II698);
  IV  NOT_297(II709,n275gat);
  IV  NOT_298(n274gat,II709);
  IV  NOT_299(II712,n274gat);
  IV  NOT_300(n348gat,II712);
  IV  NOT_301(II715,n401gat);
  IV  NOT_302(n349gat,II715);
  IV  NOT_303(II718,n398gat);
  IV  NOT_304(n397gat,II718);
  IV  NOT_305(II721,n397gat);
  IV  NOT_306(n350gat,II721);
  IV  NOT_307(n400gat,n402gat);
  IV  NOT_308(II726,n400gat);
  IV  NOT_309(n351gat,II726);
  IV  NOT_310(II729,n396gat);
  IV  NOT_311(n352gat,II729);
  IV  NOT_312(n273gat,n275gat);
  IV  NOT_313(II734,n273gat);
  IV  NOT_314(n353gat,II734);
  IV  NOT_315(n178gat,n343gat);
  IV  NOT_316(II741,n178gat);
  IV  NOT_317(n62gat,II741);
  IV  NOT_318(n66gat,n906gat);
  IV  NOT_319(II746,n66gat);
  IV  NOT_320(n63gat,II746);
  IV  NOT_321(II749,n343gat);
  IV  NOT_322(n64gat,II749);
  IV  NOT_323(II753,n167gat);
  IV  NOT_324(n65gat,II753);
  IV  NOT_325(n2474gat,n2476gat);
  IV  NOT_326(II768,n3090gat);
  IV  NOT_327(n2832gat,II768);
  IV  NOT_328(II771,n2832gat);
  IV  NOT_329(n2831gat,II771);
  IV  NOT_330(n2731gat,n2733gat);
  IV  NOT_331(II776,n3074gat);
  IV  NOT_332(n2719gat,II776);
  IV  NOT_333(n2718gat,n2719gat);
  IV  NOT_334(II790,n1068gat);
  IV  NOT_335(n1067gat,II790);
  IV  NOT_336(II793,n1067gat);
  IV  NOT_337(n949gat,II793);
  IV  NOT_338(II796,n3076gat);
  IV  NOT_339(n2839gat,II796);
  IV  NOT_340(n2838gat,n2839gat);
  IV  NOT_341(n2775gat,n2777gat);
  IV  NOT_342(II812,n957gat);
  IV  NOT_343(n956gat,II812);
  IV  NOT_344(II815,n956gat);
  IV  NOT_345(n950gat,II815);
  IV  NOT_346(II818,n3075gat);
  IV  NOT_347(n2712gat,II818);
  IV  NOT_348(n2711gat,n2712gat);
  IV  NOT_349(n2734gat,n2736gat);
  IV  NOT_350(II834,n861gat);
  IV  NOT_351(n860gat,II834);
  IV  NOT_352(II837,n860gat);
  IV  NOT_353(n951gat,II837);
  IV  NOT_354(n955gat,n957gat);
  IV  NOT_355(II842,n955gat);
  IV  NOT_356(n952gat,II842);
  IV  NOT_357(n859gat,n861gat);
  IV  NOT_358(II846,n859gat);
  IV  NOT_359(n953gat,II846);
  IV  NOT_360(n1066gat,n1068gat);
  IV  NOT_361(II851,n1066gat);
  IV  NOT_362(n954gat,II851);
  IV  NOT_363(n857gat,n944gat);
  IV  NOT_364(II858,n857gat);
  IV  NOT_365(n938gat,II858);
  IV  NOT_366(n2792gat,n2794gat);
  IV  NOT_367(II863,n3080gat);
  IV  NOT_368(n2847gat,II863);
  IV  NOT_369(n2846gat,n2847gat);
  IV  NOT_370(II877,n1294gat);
  IV  NOT_371(n1293gat,II877);
  IV  NOT_372(II880,n1293gat);
  IV  NOT_373(n1233gat,II880);
  IV  NOT_374(n2672gat,n2674gat);
  IV  NOT_375(II885,n3082gat);
  IV  NOT_376(n2853gat,II885);
  IV  NOT_377(n2852gat,n2853gat);
  IV  NOT_378(II899,n1241gat);
  IV  NOT_379(n1240gat,II899);
  IV  NOT_380(II902,n1240gat);
  IV  NOT_381(n1234gat,II902);
  IV  NOT_382(II913,n1298gat);
  IV  NOT_383(n1297gat,II913);
  IV  NOT_384(II916,n1297gat);
  IV  NOT_385(n1235gat,II916);
  IV  NOT_386(n1239gat,n1241gat);
  IV  NOT_387(II921,n1239gat);
  IV  NOT_388(n1236gat,II921);
  IV  NOT_389(n1296gat,n1298gat);
  IV  NOT_390(II925,n1296gat);
  IV  NOT_391(n1237gat,II925);
  IV  NOT_392(n1292gat,n1294gat);
  IV  NOT_393(II930,n1292gat);
  IV  NOT_394(n1238gat,II930);
  IV  NOT_395(II936,n1228gat);
  IV  NOT_396(n939gat,II936);
  IV  NOT_397(n2778gat,n2780gat);
  IV  NOT_398(II941,n3077gat);
  IV  NOT_399(n2837gat,II941);
  IV  NOT_400(n2836gat,n2837gat);
  IV  NOT_401(II955,n865gat);
  IV  NOT_402(n864gat,II955);
  IV  NOT_403(II958,n864gat);
  IV  NOT_404(n1055gat,II958);
  IV  NOT_405(n2789gat,n2791gat);
  IV  NOT_406(II963,n3079gat);
  IV  NOT_407(n2841gat,II963);
  IV  NOT_408(n2840gat,n2841gat);
  IV  NOT_409(II977,n1080gat);
  IV  NOT_410(n1079gat,II977);
  IV  NOT_411(II980,n1079gat);
  IV  NOT_412(n1056gat,II980);
  IV  NOT_413(n2781gat,n2783gat);
  IV  NOT_414(II985,n3078gat);
  IV  NOT_415(n2843gat,II985);
  IV  NOT_416(n2842gat,n2843gat);
  IV  NOT_417(II999,n1148gat);
  IV  NOT_418(n1147gat,II999);
  IV  NOT_419(II1002,n1147gat);
  IV  NOT_420(n1057gat,II1002);
  IV  NOT_421(n1078gat,n1080gat);
  IV  NOT_422(II1007,n1078gat);
  IV  NOT_423(n1058gat,II1007);
  IV  NOT_424(n1146gat,n1148gat);
  IV  NOT_425(II1011,n1146gat);
  IV  NOT_426(n1059gat,II1011);
  IV  NOT_427(n863gat,n865gat);
  IV  NOT_428(II1016,n863gat);
  IV  NOT_429(n1060gat,II1016);
  IV  NOT_430(n928gat,n1050gat);
  IV  NOT_431(II1023,n928gat);
  IV  NOT_432(n940gat,II1023);
  IV  NOT_433(n858gat,n1228gat);
  IV  NOT_434(II1028,n858gat);
  IV  NOT_435(n941gat,II1028);
  IV  NOT_436(II1031,n1050gat);
  IV  NOT_437(n942gat,II1031);
  IV  NOT_438(II1035,n944gat);
  IV  NOT_439(n943gat,II1035);
  IV  NOT_440(n2466gat,n2468gat);
  IV  NOT_441(n2720gat,n2722gat);
  IV  NOT_442(n740gat,n2667gat);
  IV  NOT_443(n2784gat,n2786gat);
  IV  NOT_444(n743gat,n746gat);
  IV  NOT_445(n294gat,n360gat);
  IV  NOT_446(n374gat,n2767gat);
  IV  NOT_447(n616gat,n618gat);
  IV  NOT_448(II1067,n616gat);
  IV  NOT_449(n501gat,II1067);
  IV  NOT_450(n489gat,n491gat);
  IV  NOT_451(II1079,n489gat);
  IV  NOT_452(n502gat,II1079);
  IV  NOT_453(II1082,n618gat);
  IV  NOT_454(n617gat,II1082);
  IV  NOT_455(II1085,n617gat);
  IV  NOT_456(n499gat,II1085);
  IV  NOT_457(II1088,n491gat);
  IV  NOT_458(n490gat,II1088);
  IV  NOT_459(II1091,n490gat);
  IV  NOT_460(n500gat,II1091);
  IV  NOT_461(n620gat,n622gat);
  IV  NOT_462(II1103,n620gat);
  IV  NOT_463(n738gat,II1103);
  IV  NOT_464(n624gat,n626gat);
  IV  NOT_465(II1115,n624gat);
  IV  NOT_466(n737gat,II1115);
  IV  NOT_467(II1118,n622gat);
  IV  NOT_468(n621gat,II1118);
  IV  NOT_469(II1121,n621gat);
  IV  NOT_470(n733gat,II1121);
  IV  NOT_471(II1124,n626gat);
  IV  NOT_472(n625gat,II1124);
  IV  NOT_473(II1127,n625gat);
  IV  NOT_474(n735gat,II1127);
  IV  NOT_475(II1138,n834gat);
  IV  NOT_476(n833gat,II1138);
  IV  NOT_477(II1141,n833gat);
  IV  NOT_478(n714gat,II1141);
  IV  NOT_479(II1152,n707gat);
  IV  NOT_480(n706gat,II1152);
  IV  NOT_481(II1155,n706gat);
  IV  NOT_482(n715gat,II1155);
  IV  NOT_483(II1166,n838gat);
  IV  NOT_484(n837gat,II1166);
  IV  NOT_485(II1169,n837gat);
  IV  NOT_486(n716gat,II1169);
  IV  NOT_487(n705gat,n707gat);
  IV  NOT_488(II1174,n705gat);
  IV  NOT_489(n717gat,II1174);
  IV  NOT_490(n836gat,n838gat);
  IV  NOT_491(II1178,n836gat);
  IV  NOT_492(n718gat,II1178);
  IV  NOT_493(n832gat,n834gat);
  IV  NOT_494(II1183,n832gat);
  IV  NOT_495(n719gat,II1183);
  IV  NOT_496(n515gat,n709gat);
  IV  NOT_497(II1190,n515gat);
  IV  NOT_498(n509gat,II1190);
  IV  NOT_499(II1201,n830gat);
  IV  NOT_500(n829gat,II1201);
  IV  NOT_501(II1204,n829gat);
  IV  NOT_502(n734gat,II1204);
  IV  NOT_503(n828gat,n830gat);
  IV  NOT_504(II1209,n828gat);
  IV  NOT_505(n736gat,II1209);
  IV  NOT_506(II1216,n728gat);
  IV  NOT_507(n510gat,II1216);
  IV  NOT_508(II1227,n614gat);
  IV  NOT_509(n613gat,II1227);
  IV  NOT_510(II1230,n613gat);
  IV  NOT_511(n498gat,II1230);
  IV  NOT_512(n612gat,n614gat);
  IV  NOT_513(II1236,n612gat);
  IV  NOT_514(n503gat,II1236);
  IV  NOT_515(n404gat,n493gat);
  IV  NOT_516(II1243,n404gat);
  IV  NOT_517(n511gat,II1243);
  IV  NOT_518(n405gat,n728gat);
  IV  NOT_519(II1248,n405gat);
  IV  NOT_520(n512gat,II1248);
  IV  NOT_521(II1251,n493gat);
  IV  NOT_522(n513gat,II1251);
  IV  NOT_523(II1255,n709gat);
  IV  NOT_524(n514gat,II1255);
  IV  NOT_525(n2524gat,n2526gat);
  IV  NOT_526(n17gat,n564gat);
  IV  NOT_527(n79gat,n86gat);
  IV  NOT_528(n219gat,n78gat);
  IV  NOT_529(n563gat,II1278);
  IV  NOT_530(n289gat,n563gat);
  IV  NOT_531(n179gat,n287gat);
  IV  NOT_532(n188gat,n288gat);
  IV  NOT_533(n72gat,n181gat);
  IV  NOT_534(n111gat,n182gat);
  IV  NOT_535(II1302,n680gat);
  IV  NOT_536(n679gat,II1302);
  IV  NOT_537(II1305,n679gat);
  IV  NOT_538(n808gat,II1305);
  IV  NOT_539(II1319,n816gat);
  IV  NOT_540(n815gat,II1319);
  IV  NOT_541(II1322,n815gat);
  IV  NOT_542(n809gat,II1322);
  IV  NOT_543(II1336,n580gat);
  IV  NOT_544(n579gat,II1336);
  IV  NOT_545(II1339,n579gat);
  IV  NOT_546(n810gat,II1339);
  IV  NOT_547(n814gat,n816gat);
  IV  NOT_548(II1344,n814gat);
  IV  NOT_549(n811gat,II1344);
  IV  NOT_550(n578gat,n580gat);
  IV  NOT_551(II1348,n578gat);
  IV  NOT_552(n812gat,II1348);
  IV  NOT_553(n678gat,n680gat);
  IV  NOT_554(II1353,n678gat);
  IV  NOT_555(n813gat,II1353);
  IV  NOT_556(n677gat,n803gat);
  IV  NOT_557(II1360,n677gat);
  IV  NOT_558(n572gat,II1360);
  IV  NOT_559(II1371,n824gat);
  IV  NOT_560(n823gat,II1371);
  IV  NOT_561(II1374,n823gat);
  IV  NOT_562(n591gat,II1374);
  IV  NOT_563(II1385,n820gat);
  IV  NOT_564(n819gat,II1385);
  IV  NOT_565(II1388,n819gat);
  IV  NOT_566(n592gat,II1388);
  IV  NOT_567(II1399,n883gat);
  IV  NOT_568(n882gat,II1399);
  IV  NOT_569(II1402,n882gat);
  IV  NOT_570(n593gat,II1402);
  IV  NOT_571(n818gat,n820gat);
  IV  NOT_572(II1407,n818gat);
  IV  NOT_573(n594gat,II1407);
  IV  NOT_574(n881gat,n883gat);
  IV  NOT_575(II1411,n881gat);
  IV  NOT_576(n595gat,II1411);
  IV  NOT_577(n822gat,n824gat);
  IV  NOT_578(II1416,n822gat);
  IV  NOT_579(n596gat,II1416);
  IV  NOT_580(II1422,n586gat);
  IV  NOT_581(n573gat,II1422);
  IV  NOT_582(II1436,n584gat);
  IV  NOT_583(n583gat,II1436);
  IV  NOT_584(II1439,n583gat);
  IV  NOT_585(n691gat,II1439);
  IV  NOT_586(II1450,n684gat);
  IV  NOT_587(n683gat,II1450);
  IV  NOT_588(II1453,n683gat);
  IV  NOT_589(n692gat,II1453);
  IV  NOT_590(II1464,n699gat);
  IV  NOT_591(n698gat,II1464);
  IV  NOT_592(II1467,n698gat);
  IV  NOT_593(n693gat,II1467);
  IV  NOT_594(n682gat,n684gat);
  IV  NOT_595(II1472,n682gat);
  IV  NOT_596(n694gat,II1472);
  IV  NOT_597(n697gat,n699gat);
  IV  NOT_598(II1476,n697gat);
  IV  NOT_599(n695gat,II1476);
  IV  NOT_600(n582gat,n584gat);
  IV  NOT_601(II1481,n582gat);
  IV  NOT_602(n696gat,II1481);
  IV  NOT_603(n456gat,n686gat);
  IV  NOT_604(II1488,n456gat);
  IV  NOT_605(n574gat,II1488);
  IV  NOT_606(n565gat,n586gat);
  IV  NOT_607(II1493,n565gat);
  IV  NOT_608(n575gat,II1493);
  IV  NOT_609(II1496,n686gat);
  IV  NOT_610(n576gat,II1496);
  IV  NOT_611(II1500,n803gat);
  IV  NOT_612(n577gat,II1500);
  IV  NOT_613(n2462gat,n2464gat);
  IV  NOT_614(n2665gat,II1516);
  IV  NOT_615(n2596gat,n2665gat);
  IV  NOT_616(n189gat,n286gat);
  IV  NOT_617(n194gat,n187gat);
  IV  NOT_618(n21gat,n15gat);
  IV  NOT_619(II1538,n2399gat);
  IV  NOT_620(n2398gat,II1538);
  IV  NOT_621(n2353gat,n2398gat);
  IV  NOT_622(II1550,n2343gat);
  IV  NOT_623(n2342gat,II1550);
  IV  NOT_624(n2284gat,n2342gat);
  IV  NOT_625(n2201gat,n2203gat);
  IV  NOT_626(n2354gat,n2201gat);
  IV  NOT_627(n2560gat,n2562gat);
  IV  NOT_628(n2356gat,n2560gat);
  IV  NOT_629(n2205gat,n2207gat);
  IV  NOT_630(n2214gat,n2205gat);
  IV  NOT_631(n2286gat,II1585);
  IV  NOT_632(n2624gat,n2626gat);
  IV  NOT_633(II1606,n2490gat);
  IV  NOT_634(n2489gat,II1606);
  IV  NOT_635(II1617,n2622gat);
  IV  NOT_636(n2621gat,II1617);
  IV  NOT_637(n2533gat,n2534gat);
  IV  NOT_638(II1630,n2630gat);
  IV  NOT_639(n2629gat,II1630);
  IV  NOT_640(n2486gat,n2629gat);
  IV  NOT_641(n2541gat,n2543gat);
  IV  NOT_642(n2429gat,n2541gat);
  IV  NOT_643(n2432gat,n2430gat);
  IV  NOT_644(II1655,n2102gat);
  IV  NOT_645(n2101gat,II1655);
  IV  NOT_646(n1693gat,n2101gat);
  IV  NOT_647(II1667,n1880gat);
  IV  NOT_648(n1879gat,II1667);
  IV  NOT_649(n1698gat,n1934gat);
  IV  NOT_650(n1543gat,n1606gat);
  IV  NOT_651(II1683,n1763gat);
  IV  NOT_652(n1762gat,II1683);
  IV  NOT_653(n1673gat,n2989gat);
  IV  NOT_654(n1858gat,n1673gat);
  IV  NOT_655(II1698,n2155gat);
  IV  NOT_656(n2154gat,II1698);
  IV  NOT_657(n2488gat,n2490gat);
  IV  NOT_658(II1703,n2626gat);
  IV  NOT_659(n2625gat,II1703);
  IV  NOT_660(n2530gat,n2531gat);
  IV  NOT_661(II1708,n2543gat);
  IV  NOT_662(n2542gat,II1708);
  IV  NOT_663(n2482gat,n2542gat);
  IV  NOT_664(n2426gat,n2480gat);
  IV  NOT_665(n2153gat,n2155gat);
  IV  NOT_666(n2341gat,n2343gat);
  IV  NOT_667(n2355gat,n2341gat);
  IV  NOT_668(II1719,n2562gat);
  IV  NOT_669(n2561gat,II1719);
  IV  NOT_670(n2443gat,n2561gat);
  IV  NOT_671(n2289gat,II1724);
  IV  NOT_672(n2148gat,II1734);
  IV  NOT_673(n855gat,n2148gat);
  IV  NOT_674(n759gat,n855gat);
  IV  NOT_675(II1749,n1035gat);
  IV  NOT_676(n1034gat,II1749);
  IV  NOT_677(II1752,n1034gat);
  IV  NOT_678(n1189gat,II1752);
  IV  NOT_679(n1075gat,n855gat);
  IV  NOT_680(II1766,n1121gat);
  IV  NOT_681(n1120gat,II1766);
  IV  NOT_682(II1769,n1120gat);
  IV  NOT_683(n1190gat,II1769);
  IV  NOT_684(n760gat,n855gat);
  IV  NOT_685(II1783,n1072gat);
  IV  NOT_686(n1071gat,II1783);
  IV  NOT_687(II1786,n1071gat);
  IV  NOT_688(n1191gat,II1786);
  IV  NOT_689(n1119gat,n1121gat);
  IV  NOT_690(II1791,n1119gat);
  IV  NOT_691(n1192gat,II1791);
  IV  NOT_692(n1070gat,n1072gat);
  IV  NOT_693(II1795,n1070gat);
  IV  NOT_694(n1193gat,II1795);
  IV  NOT_695(n1033gat,n1035gat);
  IV  NOT_696(II1800,n1033gat);
  IV  NOT_697(n1194gat,II1800);
  IV  NOT_698(n1183gat,n1184gat);
  IV  NOT_699(II1807,n1183gat);
  IV  NOT_700(n1274gat,II1807);
  IV  NOT_701(n644gat,n855gat);
  IV  NOT_702(n1280gat,n1282gat);
  IV  NOT_703(n641gat,n855gat);
  IV  NOT_704(II1833,n1226gat);
  IV  NOT_705(n1225gat,II1833);
  IV  NOT_706(II1837,n1282gat);
  IV  NOT_707(n1281gat,II1837);
  IV  NOT_708(n1224gat,n1226gat);
  IV  NOT_709(II1843,n2970gat);
  IV  NOT_710(n1275gat,II1843);
  IV  NOT_711(n761gat,n855gat);
  IV  NOT_712(II1857,n931gat);
  IV  NOT_713(n930gat,II1857);
  IV  NOT_714(II1860,n930gat);
  IV  NOT_715(n1206gat,II1860);
  IV  NOT_716(n762gat,n855gat);
  IV  NOT_717(II1874,n1135gat);
  IV  NOT_718(n1134gat,II1874);
  IV  NOT_719(II1877,n1134gat);
  IV  NOT_720(n1207gat,II1877);
  IV  NOT_721(n643gat,n855gat);
  IV  NOT_722(II1891,n1045gat);
  IV  NOT_723(n1044gat,II1891);
  IV  NOT_724(II1894,n1044gat);
  IV  NOT_725(n1208gat,II1894);
  IV  NOT_726(n1133gat,n1135gat);
  IV  NOT_727(II1899,n1133gat);
  IV  NOT_728(n1209gat,II1899);
  IV  NOT_729(n1043gat,n1045gat);
  IV  NOT_730(II1903,n1043gat);
  IV  NOT_731(n1210gat,II1903);
  IV  NOT_732(n929gat,n931gat);
  IV  NOT_733(II1908,n929gat);
  IV  NOT_734(n1211gat,II1908);
  IV  NOT_735(n1268gat,n1201gat);
  IV  NOT_736(II1915,n1268gat);
  IV  NOT_737(n1276gat,II1915);
  IV  NOT_738(n1329gat,n2970gat);
  IV  NOT_739(II1920,n1329gat);
  IV  NOT_740(n1277gat,II1920);
  IV  NOT_741(II1923,n1201gat);
  IV  NOT_742(n1278gat,II1923);
  IV  NOT_743(II1927,n1184gat);
  IV  NOT_744(n1279gat,II1927);
  IV  NOT_745(n1284gat,n1269gat);
  IV  NOT_746(n642gat,n855gat);
  IV  NOT_747(n1195gat,n1197gat);
  IV  NOT_748(II1947,n1197gat);
  IV  NOT_749(n1196gat,II1947);
  IV  NOT_750(n2516gat,n2518gat);
  IV  NOT_751(II1961,n2516gat);
  IV  NOT_752(n3017gat,II1961);
  IV  NOT_753(n851gat,n853gat);
  IV  NOT_754(n1725gat,n2148gat);
  IV  NOT_755(n664gat,n1725gat);
  IV  NOT_756(n852gat,n854gat);
  IV  NOT_757(II1981,n667gat);
  IV  NOT_758(n666gat,II1981);
  IV  NOT_759(n368gat,n1725gat);
  IV  NOT_760(II1996,n659gat);
  IV  NOT_761(n658gat,II1996);
  IV  NOT_762(II1999,n658gat);
  IV  NOT_763(n784gat,II1999);
  IV  NOT_764(n662gat,n1725gat);
  IV  NOT_765(II2014,n553gat);
  IV  NOT_766(n552gat,II2014);
  IV  NOT_767(II2017,n552gat);
  IV  NOT_768(n785gat,II2017);
  IV  NOT_769(n661gat,n1725gat);
  IV  NOT_770(II2032,n777gat);
  IV  NOT_771(n776gat,II2032);
  IV  NOT_772(II2035,n776gat);
  IV  NOT_773(n786gat,II2035);
  IV  NOT_774(n551gat,n553gat);
  IV  NOT_775(II2040,n551gat);
  IV  NOT_776(n787gat,II2040);
  IV  NOT_777(n775gat,n777gat);
  IV  NOT_778(II2044,n775gat);
  IV  NOT_779(n788gat,II2044);
  IV  NOT_780(n657gat,n659gat);
  IV  NOT_781(II2049,n657gat);
  IV  NOT_782(n789gat,II2049);
  IV  NOT_783(n35gat,n779gat);
  IV  NOT_784(II2056,n35gat);
  IV  NOT_785(n125gat,II2056);
  IV  NOT_786(n558gat,n1725gat);
  IV  NOT_787(n559gat,n561gat);
  IV  NOT_788(n371gat,n1725gat);
  IV  NOT_789(II2084,n366gat);
  IV  NOT_790(n365gat,II2084);
  IV  NOT_791(II2088,n561gat);
  IV  NOT_792(n560gat,II2088);
  IV  NOT_793(n364gat,n366gat);
  IV  NOT_794(II2094,n2876gat);
  IV  NOT_795(n126gat,II2094);
  IV  NOT_796(n663gat,n1725gat);
  IV  NOT_797(II2109,n322gat);
  IV  NOT_798(n321gat,II2109);
  IV  NOT_799(II2112,n321gat);
  IV  NOT_800(n226gat,II2112);
  IV  NOT_801(n370gat,n1725gat);
  IV  NOT_802(II2127,n318gat);
  IV  NOT_803(n317gat,II2127);
  IV  NOT_804(II2130,n317gat);
  IV  NOT_805(n227gat,II2130);
  IV  NOT_806(n369gat,n1725gat);
  IV  NOT_807(II2145,n314gat);
  IV  NOT_808(n313gat,II2145);
  IV  NOT_809(II2148,n313gat);
  IV  NOT_810(n228gat,II2148);
  IV  NOT_811(n316gat,n318gat);
  IV  NOT_812(II2153,n316gat);
  IV  NOT_813(n229gat,II2153);
  IV  NOT_814(n312gat,n314gat);
  IV  NOT_815(II2157,n312gat);
  IV  NOT_816(n230gat,II2157);
  IV  NOT_817(n320gat,n322gat);
  IV  NOT_818(II2162,n320gat);
  IV  NOT_819(n231gat,II2162);
  IV  NOT_820(n34gat,n221gat);
  IV  NOT_821(II2169,n34gat);
  IV  NOT_822(n127gat,II2169);
  IV  NOT_823(n133gat,n2876gat);
  IV  NOT_824(II2174,n133gat);
  IV  NOT_825(n128gat,II2174);
  IV  NOT_826(II2177,n221gat);
  IV  NOT_827(n129gat,II2177);
  IV  NOT_828(II2181,n779gat);
  IV  NOT_829(n130gat,II2181);
  IV  NOT_830(n665gat,n667gat);
  IV  NOT_831(n1601gat,n120gat);
  IV  NOT_832(n2597gat,n2599gat);
  IV  NOT_833(n2595gat,n2594gat);
  IV  NOT_834(n2586gat,n2588gat);
  IV  NOT_835(II2213,n2342gat);
  IV  NOT_836(n2573gat,II2213);
  IV  NOT_837(n2638gat,n2640gat);
  IV  NOT_838(II2225,n2638gat);
  IV  NOT_839(n2574gat,II2225);
  IV  NOT_840(II2228,n2561gat);
  IV  NOT_841(n2575gat,II2228);
  IV  NOT_842(II2232,n2640gat);
  IV  NOT_843(n2639gat,II2232);
  IV  NOT_844(II2235,n2639gat);
  IV  NOT_845(n2576gat,II2235);
  IV  NOT_846(II2238,n2560gat);
  IV  NOT_847(n2577gat,II2238);
  IV  NOT_848(II2242,n2341gat);
  IV  NOT_849(n2578gat,II2242);
  IV  NOT_850(II2248,n2568gat);
  IV  NOT_851(n2582gat,II2248);
  IV  NOT_852(II2251,n2207gat);
  IV  NOT_853(n2206gat,II2251);
  IV  NOT_854(II2254,n2206gat);
  IV  NOT_855(n2414gat,II2254);
  IV  NOT_856(II2257,n2398gat);
  IV  NOT_857(n2415gat,II2257);
  IV  NOT_858(II2260,n2203gat);
  IV  NOT_859(n2202gat,II2260);
  IV  NOT_860(II2263,n2202gat);
  IV  NOT_861(n2416gat,II2263);
  IV  NOT_862(n2397gat,n2399gat);
  IV  NOT_863(II2268,n2397gat);
  IV  NOT_864(n2417gat,II2268);
  IV  NOT_865(II2271,n2201gat);
  IV  NOT_866(n2418gat,II2271);
  IV  NOT_867(II2275,n2205gat);
  IV  NOT_868(n2419gat,II2275);
  IV  NOT_869(II2281,n2409gat);
  IV  NOT_870(n2585gat,II2281);
  IV  NOT_871(n2656gat,n2658gat);
  IV  NOT_872(n2493gat,n2495gat);
  IV  NOT_873(n2388gat,n2390gat);
  IV  NOT_874(II2316,n2390gat);
  IV  NOT_875(n2389gat,II2316);
  IV  NOT_876(II2319,n2495gat);
  IV  NOT_877(n2494gat,II2319);
  IV  NOT_878(II2324,n3014gat);
  IV  NOT_879(n2649gat,II2324);
  IV  NOT_880(n2268gat,n2270gat);
  IV  NOT_881(II2344,n2339gat);
  IV  NOT_882(n2338gat,II2344);
  IV  NOT_883(n2337gat,n2339gat);
  IV  NOT_884(II2349,n2270gat);
  IV  NOT_885(n2269gat,II2349);
  IV  NOT_886(II2354,n2880gat);
  IV  NOT_887(n2652gat,II2354);
  IV  NOT_888(n2500gat,n2502gat);
  IV  NOT_889(n2620gat,n2622gat);
  IV  NOT_890(n2612gat,n2620gat);
  IV  NOT_891(II2372,n2612gat);
  IV  NOT_892(n2606gat,II2372);
  IV  NOT_893(n2532gat,n2625gat);
  IV  NOT_894(II2376,n2532gat);
  IV  NOT_895(n2607gat,II2376);
  IV  NOT_896(n2540gat,n2488gat);
  IV  NOT_897(II2380,n2540gat);
  IV  NOT_898(n2608gat,II2380);
  IV  NOT_899(n2536gat,n2624gat);
  IV  NOT_900(II2385,n2536gat);
  IV  NOT_901(n2609gat,II2385);
  IV  NOT_902(n2487gat,n2489gat);
  IV  NOT_903(II2389,n2487gat);
  IV  NOT_904(n2610gat,II2389);
  IV  NOT_905(n2557gat,n2621gat);
  IV  NOT_906(II2394,n2557gat);
  IV  NOT_907(n2611gat,II2394);
  IV  NOT_908(II2400,n2601gat);
  IV  NOT_909(n2616gat,II2400);
  IV  NOT_910(II2403,n2629gat);
  IV  NOT_911(n2550gat,II2403);
  IV  NOT_912(II2414,n2634gat);
  IV  NOT_913(n2633gat,II2414);
  IV  NOT_914(II2417,n2633gat);
  IV  NOT_915(n2551gat,II2417);
  IV  NOT_916(II2420,n2542gat);
  IV  NOT_917(n2552gat,II2420);
  IV  NOT_918(n2632gat,n2634gat);
  IV  NOT_919(II2425,n2632gat);
  IV  NOT_920(n2553gat,II2425);
  IV  NOT_921(II2428,n2541gat);
  IV  NOT_922(n2554gat,II2428);
  IV  NOT_923(n2628gat,n2630gat);
  IV  NOT_924(II2433,n2628gat);
  IV  NOT_925(n2555gat,II2433);
  IV  NOT_926(II2439,n2545gat);
  IV  NOT_927(n2619gat,II2439);
  IV  NOT_928(n2504gat,n2506gat);
  IV  NOT_929(n2660gat,n2655gat);
  IV  NOT_930(n1528gat,n2293gat);
  IV  NOT_931(n1523gat,n2219gat);
  IV  NOT_932(n1592gat,n1529gat);
  IV  NOT_933(n2666gat,n1704gat);
  IV  NOT_934(n2422gat,n3013gat);
  IV  NOT_935(n2290gat,n2202gat);
  IV  NOT_936(n2081gat,n2218gat);
  IV  NOT_937(n2285gat,n2397gat);
  IV  NOT_938(n2359gat,n2358gat);
  IV  NOT_939(n1414gat,n1415gat);
  IV  NOT_940(n566gat,n364gat);
  IV  NOT_941(n1480gat,n2292gat);
  IV  NOT_942(n1301gat,n1416gat);
  IV  NOT_943(n1150gat,n312gat);
  IV  NOT_944(n873gat,n316gat);
  IV  NOT_945(n2011gat,n2306gat);
  IV  NOT_946(n1478gat,n1481gat);
  IV  NOT_947(n875gat,n559gat);
  IV  NOT_948(n1410gat,n2357gat);
  IV  NOT_949(n876gat,n1347gat);
  IV  NOT_950(n1160gat,n1484gat);
  IV  NOT_951(n1084gat,n657gat);
  IV  NOT_952(n983gat,n320gat);
  IV  NOT_953(n1482gat,n2363gat);
  IV  NOT_954(n1157gat,n1483gat);
  IV  NOT_955(n985gat,n775gat);
  IV  NOT_956(n1530gat,n2364gat);
  IV  NOT_957(n1307gat,n1308gat);
  IV  NOT_958(n1085gat,n551gat);
  IV  NOT_959(n1479gat,n2291gat);
  IV  NOT_960(n1348gat,n1349gat);
  IV  NOT_961(n2217gat,n2206gat);
  IV  NOT_962(n1591gat,n2223gat);
  IV  NOT_963(n1437gat,n1438gat);
  IV  NOT_964(n1832gat,n1834gat);
  IV  NOT_965(n1765gat,n1767gat);
  IV  NOT_966(n1878gat,n1880gat);
  IV  NOT_967(n1442gat,n1831gat);
  IV  NOT_968(n1444gat,n1442gat);
  IV  NOT_969(n1378gat,n2975gat);
  IV  NOT_970(n1322gat,n2974gat);
  IV  NOT_971(n1439gat,n1486gat);
  IV  NOT_972(n1370gat,n1426gat);
  IV  NOT_973(n1369gat,n2966gat);
  IV  NOT_974(n1366gat,n1365gat);
  IV  NOT_975(n1374gat,n2979gat);
  IV  NOT_976(n2162gat,n2220gat);
  IV  NOT_977(n1450gat,n1423gat);
  IV  NOT_978(n1427gat,n1608gat);
  IV  NOT_979(n1603gat,n1831gat);
  IV  NOT_980(n2082gat,n2084gat);
  IV  NOT_981(n1449gat,n1494gat);
  IV  NOT_982(n1590gat,n1603gat);
  IV  NOT_983(n1248gat,n2954gat);
  IV  NOT_984(n1418gat,n1417gat);
  IV  NOT_985(n1306gat,n2964gat);
  IV  NOT_986(n1353gat,n1419gat);
  IV  NOT_987(n1247gat,n2958gat);
  IV  NOT_988(n1355gat,n1422gat);
  IV  NOT_989(n1300gat,n2963gat);
  IV  NOT_990(n1487gat,n1485gat);
  IV  NOT_991(n1164gat,n2953gat);
  IV  NOT_992(n1356gat,n1354gat);
  IV  NOT_993(n1436gat,n1435gat);
  IV  NOT_994(n1106gat,n2949gat);
  IV  NOT_995(n1425gat,n1421gat);
  IV  NOT_996(n1105gat,n2934gat);
  IV  NOT_997(n1424gat,n1420gat);
  IV  NOT_998(n1309gat,n2959gat);
  IV  NOT_999(II2672,n2143gat);
  IV  NOT_1000(n2142gat,II2672);
  IV  NOT_1001(n1788gat,n2142gat);
  IV  NOT_1002(II2684,n2061gat);
  IV  NOT_1003(n2060gat,II2684);
  IV  NOT_1004(n1786gat,n2060gat);
  IV  NOT_1005(II2696,n2139gat);
  IV  NOT_1006(n2138gat,II2696);
  IV  NOT_1007(n1839gat,n2138gat);
  IV  NOT_1008(n1897gat,n1899gat);
  IV  NOT_1009(n1884gat,n1897gat);
  IV  NOT_1010(n1848gat,n1850gat);
  IV  NOT_1011(n1783gat,n1848gat);
  IV  NOT_1012(n1548gat,II2721);
  IV  NOT_1013(n1719gat,n1548gat);
  IV  NOT_1014(n2137gat,n2139gat);
  IV  NOT_1015(n1633gat,n2137gat);
  IV  NOT_1016(n2059gat,n2061gat);
  IV  NOT_1017(n1785gat,n2059gat);
  IV  NOT_1018(II2731,n1850gat);
  IV  NOT_1019(n1849gat,II2731);
  IV  NOT_1020(n1784gat,n1849gat);
  IV  NOT_1021(n1716gat,II2736);
  IV  NOT_1022(n1635gat,n1716gat);
  IV  NOT_1023(n2401gat,n2403gat);
  IV  NOT_1024(n1989gat,n2401gat);
  IV  NOT_1025(n2392gat,n2394gat);
  IV  NOT_1026(n1918gat,n2392gat);
  IV  NOT_1027(II2771,n2440gat);
  IV  NOT_1028(n2439gat,II2771);
  IV  NOT_1029(n1986gat,n2439gat);
  IV  NOT_1030(n1866gat,n1865gat);
  IV  NOT_1031(II2785,n2407gat);
  IV  NOT_1032(n2406gat,II2785);
  IV  NOT_1033(n2216gat,n2406gat);
  IV  NOT_1034(n2345gat,n2347gat);
  IV  NOT_1035(n1988gat,n2345gat);
  IV  NOT_1036(n1735gat,n1861gat);
  IV  NOT_1037(n1387gat,n1389gat);
  IV  NOT_1038(n1694gat,II2813);
  IV  NOT_1039(n1777gat,n1694gat);
  IV  NOT_1040(n1781gat,n1780gat);
  IV  NOT_1041(n2019gat,n2021gat);
  IV  NOT_1042(n1549gat,II2832);
  IV  NOT_1043(n1551gat,n1549gat);
  IV  NOT_1044(II2837,n2347gat);
  IV  NOT_1045(n2346gat,II2837);
  IV  NOT_1046(n2152gat,n2346gat);
  IV  NOT_1047(n2405gat,n2407gat);
  IV  NOT_1048(n2351gat,n2405gat);
  IV  NOT_1049(II2843,n2403gat);
  IV  NOT_1050(n2402gat,II2843);
  IV  NOT_1051(n2212gat,n2402gat);
  IV  NOT_1052(II2847,n2394gat);
  IV  NOT_1053(n2393gat,II2847);
  IV  NOT_1054(n1991gat,n2393gat);
  IV  NOT_1055(n1665gat,n1666gat);
  IV  NOT_1056(n1517gat,n1578gat);
  IV  NOT_1057(n1392gat,n1394gat);
  IV  NOT_1058(II2873,n1496gat);
  IV  NOT_1059(n1495gat,II2873);
  IV  NOT_1060(n1685gat,n1604gat);
  IV  NOT_1061(II2885,n2091gat);
  IV  NOT_1062(n2090gat,II2885);
  IV  NOT_1063(n1550gat,II2890);
  IV  NOT_1064(n1552gat,n1550gat);
  IV  NOT_1065(n1330gat,n1332gat);
  IV  NOT_1066(n1738gat,n1740gat);
  IV  NOT_1067(II2915,n1740gat);
  IV  NOT_1068(n1739gat,II2915);
  IV  NOT_1069(n1925gat,n1920gat);
  IV  NOT_1070(n1917gat,n1921gat);
  IV  NOT_1071(n2141gat,n2143gat);
  IV  NOT_1072(n1787gat,n2141gat);
  IV  NOT_1073(n1717gat,II2926);
  IV  NOT_1074(n1859gat,n1717gat);
  IV  NOT_1075(n1922gat,n1798gat);
  IV  NOT_1076(n1713gat,II2935);
  IV  NOT_1077(n1743gat,n1713gat);
  IV  NOT_1078(n1923gat,n1864gat);
  IV  NOT_1079(n1945gat,n1690gat);
  IV  NOT_1080(II2953,n2179gat);
  IV  NOT_1081(n2178gat,II2953);
  IV  NOT_1082(n1661gat,n1660gat);
  IV  NOT_1083(n1572gat,n1576gat);
  IV  NOT_1084(n2438gat,n2440gat);
  IV  NOT_1085(n2283gat,n2438gat);
  IV  NOT_1086(n1520gat,n1582gat);
  IV  NOT_1087(n1580gat,n1577gat);
  IV  NOT_1088(n1990gat,n2988gat);
  IV  NOT_1089(II2978,n2190gat);
  IV  NOT_1090(n2189gat,II2978);
  IV  NOT_1091(II2989,n2135gat);
  IV  NOT_1092(n2134gat,II2989);
  IV  NOT_1093(II3000,n2262gat);
  IV  NOT_1094(n2261gat,II3000);
  IV  NOT_1095(n2128gat,n2129gat);
  IV  NOT_1096(n1836gat,n1695gat);
  IV  NOT_1097(II3016,n2182gat);
  IV  NOT_1098(n2181gat,II3016);
  IV  NOT_1099(n1431gat,n1433gat);
  IV  NOT_1100(n1314gat,n1316gat);
  IV  NOT_1101(n1361gat,n1363gat);
  IV  NOT_1102(II3056,n1312gat);
  IV  NOT_1103(n1311gat,II3056);
  IV  NOT_1104(n1707gat,n1626gat);
  IV  NOT_1105(n1773gat,n1775gat);
  IV  NOT_1106(n1659gat,n2987gat);
  IV  NOT_1107(n1515gat,n1521gat);
  IV  NOT_1108(n1736gat,n1737gat);
  IV  NOT_1109(n1658gat,n2216gat);
  IV  NOT_1110(n1724gat,n1732gat);
  IV  NOT_1111(n1662gat,n1663gat);
  IV  NOT_1112(n1656gat,n1655gat);
  IV  NOT_1113(n1670gat,n1667gat);
  IV  NOT_1114(n1569gat,n1570gat);
  IV  NOT_1115(n1568gat,n1575gat);
  IV  NOT_1116(n1727gat,n1728gat);
  IV  NOT_1117(n1797gat,n1801gat);
  IV  NOT_1118(n1730gat,n1731gat);
  IV  NOT_1119(n1561gat,n1571gat);
  IV  NOT_1120(n1668gat,n1734gat);
  IV  NOT_1121(n1742gat,n2216gat);
  IV  NOT_1122(n1671gat,n1669gat);
  IV  NOT_1123(n1652gat,n1657gat);
  IV  NOT_1124(n1648gat,n1729gat);
  IV  NOT_1125(n1790gat,n1726gat);
  IV  NOT_1126(n2004gat,n1929gat);
  IV  NOT_1127(n1869gat,n1871gat);
  IV  NOT_1128(II3143,n2592gat);
  IV  NOT_1129(n2591gat,II3143);
  IV  NOT_1130(n1584gat,n2989gat);
  IV  NOT_1131(n1714gat,II3149);
  IV  NOT_1132(n1718gat,n1714gat);
  IV  NOT_1133(II3163,n1508gat);
  IV  NOT_1134(n1507gat,II3163);
  IV  NOT_1135(n1396gat,n1401gat);
  IV  NOT_1136(II3168,n1394gat);
  IV  NOT_1137(n1393gat,II3168);
  IV  NOT_1138(n1409gat,n1476gat);
  IV  NOT_1139(II3174,n1899gat);
  IV  NOT_1140(n1898gat,II3174);
  IV  NOT_1141(n1838gat,n1898gat);
  IV  NOT_1142(n1712gat,II3179);
  IV  NOT_1143(II3191,n1678gat);
  IV  NOT_1144(n1677gat,II3191);
  IV  NOT_1145(n2000gat,n1412gat);
  IV  NOT_1146(n2001gat,n1412gat);
  IV  NOT_1147(n1999gat,n2001gat);
  IV  NOT_1148(n2307gat,n2309gat);
  IV  NOT_1149(II3211,n2663gat);
  IV  NOT_1150(n3018gat,II3211);
  IV  NOT_1151(n2448gat,n2450gat);
  IV  NOT_1152(n2661gat,n2662gat);
  IV  NOT_1153(n2444gat,n2446gat);
  IV  NOT_1154(II3235,n2238gat);
  IV  NOT_1155(n3019gat,II3235);
  IV  NOT_1156(n1310gat,n1312gat);
  IV  NOT_1157(n199gat,n87gat);
  IV  NOT_1158(n195gat,n184gat);
  IV  NOT_1159(n827gat,n204gat);
  IV  NOT_1160(n2093gat,n2095gat);
  IV  NOT_1161(n2174gat,n2176gat);
  IV  NOT_1162(II3273,n2169gat);
  IV  NOT_1163(n2168gat,II3273);
  IV  NOT_1164(n2452gat,n2454gat);
  IV  NOT_1165(n1691gat,n2452gat);
  IV  NOT_1166(II3287,n1691gat);
  IV  NOT_1167(n3020gat,II3287);
  IV  NOT_1168(II3290,n1691gat);
  IV  NOT_1169(n3021gat,II3290);
  IV  NOT_1170(II3293,n1691gat);
  IV  NOT_1171(n3022gat,II3293);
  IV  NOT_1172(n1699gat,n2452gat);
  IV  NOT_1173(II3297,n1699gat);
  IV  NOT_1174(n3023gat,II3297);
  IV  NOT_1175(II3300,n1699gat);
  IV  NOT_1176(n3024gat,II3300);
  IV  NOT_1177(II3303,n1691gat);
  IV  NOT_1178(n3025gat,II3303);
  IV  NOT_1179(II3306,n1699gat);
  IV  NOT_1180(n3026gat,II3306);
  IV  NOT_1181(II3309,n1699gat);
  IV  NOT_1182(n3027gat,II3309);
  IV  NOT_1183(II3312,n1699gat);
  IV  NOT_1184(n3028gat,II3312);
  IV  NOT_1185(II3315,n1869gat);
  IV  NOT_1186(n3029gat,II3315);
  IV  NOT_1187(II3318,n1869gat);
  IV  NOT_1188(n3030gat,II3318);
  IV  NOT_1189(n2260gat,n2262gat);
  IV  NOT_1190(n2257gat,n2189gat);
  IV  NOT_1191(n2188gat,n2190gat);
  IV  NOT_1192(n2187gat,n3004gat);
  IV  NOT_1193(II3336,n2040gat);
  IV  NOT_1194(n2039gat,II3336);
  IV  NOT_1195(II3339,n1775gat);
  IV  NOT_1196(n1774gat,II3339);
  IV  NOT_1197(II3342,n1316gat);
  IV  NOT_1198(n1315gat,II3342);
  IV  NOT_1199(n2042gat,n2044gat);
  IV  NOT_1200(n2035gat,n2037gat);
  IV  NOT_1201(n2023gat,n2025gat);
  IV  NOT_1202(n2097gat,n2099gat);
  IV  NOT_1203(n1855gat,n2014gat);
  IV  NOT_1204(II3387,n2194gat);
  IV  NOT_1205(n3031gat,II3387);
  IV  NOT_1206(II3390,n2261gat);
  IV  NOT_1207(n3032gat,II3390);
  IV  NOT_1208(n2256gat,n3032gat);
  IV  NOT_1209(II3394,n2260gat);
  IV  NOT_1210(n3033gat,II3394);
  IV  NOT_1211(n2251gat,n3033gat);
  IV  NOT_1212(n2184gat,n3003gat);
  IV  NOT_1213(II3401,n2192gat);
  IV  NOT_1214(n3034gat,II3401);
  IV  NOT_1215(n2133gat,n2135gat);
  IV  NOT_1216(n2131gat,n2185gat);
  IV  NOT_1217(n2049gat,n3001gat);
  IV  NOT_1218(II3412,n2057gat);
  IV  NOT_1219(n3035gat,II3412);
  IV  NOT_1220(n2253gat,n2189gat);
  IV  NOT_1221(n2252gat,n2260gat);
  IV  NOT_1222(n2248gat,n3006gat);
  IV  NOT_1223(n2264gat,n2266gat);
  IV  NOT_1224(II3429,n2266gat);
  IV  NOT_1225(n2265gat,II3429);
  IV  NOT_1226(n2492gat,n2329gat);
  IV  NOT_1227(II3436,n2492gat);
  IV  NOT_1228(n3036gat,II3436);
  IV  NOT_1229(n1709gat,n1849gat);
  IV  NOT_1230(n1845gat,n2141gat);
  IV  NOT_1231(n1891gat,n2059gat);
  IV  NOT_1232(n1963gat,n2137gat);
  IV  NOT_1233(n1886gat,n1897gat);
  IV  NOT_1234(n1968gat,n1958gat);
  IV  NOT_1235(n1629gat,n1895gat);
  IV  NOT_1236(n1631gat,n1848gat);
  IV  NOT_1237(n1711gat,n2990gat);
  IV  NOT_1238(n2200gat,n2078gat);
  IV  NOT_1239(n2437gat,n2195gat);
  IV  NOT_1240(II3457,n2556gat);
  IV  NOT_1241(n3037gat,II3457);
  IV  NOT_1242(n1956gat,n1898gat);
  IV  NOT_1243(II3461,n1956gat);
  IV  NOT_1244(n3038gat,II3461);
  IV  NOT_1245(n1954gat,n3038gat);
  IV  NOT_1246(II3465,n1886gat);
  IV  NOT_1247(n3039gat,II3465);
  IV  NOT_1248(n1888gat,n3039gat);
  IV  NOT_1249(n2048gat,n2994gat);
  IV  NOT_1250(II3472,n2539gat);
  IV  NOT_1251(n3040gat,II3472);
  IV  NOT_1252(n1969gat,n2142gat);
  IV  NOT_1253(n1893gat,n2060gat);
  IV  NOT_1254(n1892gat,n2993gat);
  IV  NOT_1255(II3483,n2436gat);
  IV  NOT_1256(n3041gat,II3483);
  IV  NOT_1257(n2056gat,n2998gat);
  IV  NOT_1258(II3491,n2387gat);
  IV  NOT_1259(n3042gat,II3491);
  IV  NOT_1260(II3494,n1963gat);
  IV  NOT_1261(n3043gat,II3494);
  IV  NOT_1262(n1960gat,n3043gat);
  IV  NOT_1263(n1887gat,n2138gat);
  IV  NOT_1264(n1961gat,n2996gat);
  IV  NOT_1265(II3504,n2330gat);
  IV  NOT_1266(n3044gat,II3504);
  IV  NOT_1267(n2199gat,n2147gat);
  IV  NOT_1268(II3509,n2438gat);
  IV  NOT_1269(n3045gat,II3509);
  IV  NOT_1270(n2332gat,n3045gat);
  IV  NOT_1271(II3513,n2439gat);
  IV  NOT_1272(n3046gat,II3513);
  IV  NOT_1273(n2259gat,n3046gat);
  IV  NOT_1274(n2328gat,n3008gat);
  IV  NOT_1275(II3520,n2498gat);
  IV  NOT_1276(n3047gat,II3520);
  IV  NOT_1277(n2151gat,n2193gat);
  IV  NOT_1278(n2209gat,n3005gat);
  IV  NOT_1279(II3530,n2396gat);
  IV  NOT_1280(n3048gat,II3530);
  IV  NOT_1281(n2052gat,n2393gat);
  IV  NOT_1282(n2058gat,n2997gat);
  IV  NOT_1283(II3539,n2198gat);
  IV  NOT_1284(n3049gat,II3539);
  IV  NOT_1285(n2349gat,n2215gat);
  IV  NOT_1286(n2281gat,n3009gat);
  IV  NOT_1287(II3549,n2197gat);
  IV  NOT_1288(n3050gat,II3549);
  IV  NOT_1289(n2146gat,n3002gat);
  IV  NOT_1290(II3558,n2196gat);
  IV  NOT_1291(n3051gat,II3558);
  IV  NOT_1292(n2031gat,n2033gat);
  IV  NOT_1293(n2108gat,n2110gat);
  IV  NOT_1294(II3587,n2125gat);
  IV  NOT_1295(n2124gat,II3587);
  IV  NOT_1296(n2123gat,n2125gat);
  IV  NOT_1297(n2119gat,n2121gat);
  IV  NOT_1298(n2115gat,n2117gat);
  IV  NOT_1299(II3610,n1882gat);
  IV  NOT_1300(n3052gat,II3610);
  IV  NOT_1301(II3621,n1975gat);
  IV  NOT_1302(n1974gat,II3621);
  IV  NOT_1303(n1955gat,n1956gat);
  IV  NOT_1304(n1970gat,n1896gat);
  IV  NOT_1305(n1973gat,n1975gat);
  IV  NOT_1306(n2558gat,n2559gat);
  IV  NOT_1307(II3635,n2558gat);
  IV  NOT_1308(n3053gat,II3635);
  IV  NOT_1309(II3646,n2644gat);
  IV  NOT_1310(n2643gat,II3646);
  IV  NOT_1311(n2333gat,n2438gat);
  IV  NOT_1312(n2564gat,n2352gat);
  IV  NOT_1313(n2642gat,n2644gat);
  IV  NOT_1314(n2636gat,n2637gat);
  IV  NOT_1315(II3660,n2636gat);
  IV  NOT_1316(n3054gat,II3660);
  IV  NOT_1317(n88gat,n84gat);
  IV  NOT_1318(n375gat,n110gat);
  IV  NOT_1319(II3677,n156gat);
  IV  NOT_1320(n155gat,II3677);
  IV  NOT_1321(n253gat,n1702gat);
  IV  NOT_1322(n150gat,n152gat);
  IV  NOT_1323(II3691,n152gat);
  IV  NOT_1324(n151gat,II3691);
  IV  NOT_1325(n243gat,n1702gat);
  IV  NOT_1326(n233gat,n243gat);
  IV  NOT_1327(n154gat,n156gat);
  IV  NOT_1328(n800gat,n2874gat);
  IV  NOT_1329(II3703,n2917gat);
  IV  NOT_1330(n3055gat,II3703);
  IV  NOT_1331(n235gat,n2878gat);
  IV  NOT_1332(II3713,n2892gat);
  IV  NOT_1333(n3056gat,II3713);
  IV  NOT_1334(n372gat,n212gat);
  IV  NOT_1335(n329gat,n331gat);
  IV  NOT_1336(II3736,n388gat);
  IV  NOT_1337(n387gat,II3736);
  IV  NOT_1338(n334gat,n1700gat);
  IV  NOT_1339(n386gat,n388gat);
  IV  NOT_1340(II3742,n331gat);
  IV  NOT_1341(n330gat,II3742);
  IV  NOT_1342(n1430gat,n1700gat);
  IV  NOT_1343(n1490gat,n1430gat);
  IV  NOT_1344(n452gat,n2885gat);
  IV  NOT_1345(II3754,n2900gat);
  IV  NOT_1346(n3057gat,II3754);
  IV  NOT_1347(n333gat,n2883gat);
  IV  NOT_1348(II3765,n2929gat);
  IV  NOT_1349(n3058gat,II3765);
  IV  NOT_1350(II3777,n463gat);
  IV  NOT_1351(n462gat,II3777);
  IV  NOT_1352(n325gat,n327gat);
  IV  NOT_1353(n457gat,n2884gat);
  IV  NOT_1354(n461gat,n463gat);
  IV  NOT_1355(n458gat,n2902gat);
  IV  NOT_1356(II3801,n2925gat);
  IV  NOT_1357(n3059gat,II3801);
  IV  NOT_1358(n144gat,n247gat);
  IV  NOT_1359(II3808,n327gat);
  IV  NOT_1360(n326gat,II3808);
  IV  NOT_1361(n878gat,n2879gat);
  IV  NOT_1362(II3817,n2916gat);
  IV  NOT_1363(n3060gat,II3817);
  IV  NOT_1364(n382gat,n384gat);
  IV  NOT_1365(II3831,n384gat);
  IV  NOT_1366(n383gat,II3831);
  IV  NOT_1367(n134gat,n2875gat);
  IV  NOT_1368(II3841,n2899gat);
  IV  NOT_1369(n3061gat,II3841);
  IV  NOT_1370(n254gat,n256gat);
  IV  NOT_1371(n252gat,n2877gat);
  IV  NOT_1372(n468gat,n470gat);
  IV  NOT_1373(II3867,n470gat);
  IV  NOT_1374(n469gat,II3867);
  IV  NOT_1375(n381gat,n2893gat);
  IV  NOT_1376(II3876,n2926gat);
  IV  NOT_1377(n3062gat,II3876);
  IV  NOT_1378(n241gat,n140gat);
  IV  NOT_1379(II3882,n256gat);
  IV  NOT_1380(n255gat,II3882);
  IV  NOT_1381(n802gat,n2882gat);
  IV  NOT_1382(II3891,n2924gat);
  IV  NOT_1383(n3063gat,II3891);
  IV  NOT_1384(n146gat,n148gat);
  IV  NOT_1385(II3904,n148gat);
  IV  NOT_1386(n147gat,II3904);
  IV  NOT_1387(n380gat,n2881gat);
  IV  NOT_1388(II3914,n2923gat);
  IV  NOT_1389(n3064gat,II3914);
  IV  NOT_1390(n69gat,n68gat);
  IV  NOT_1391(n1885gat,n2048gat);
  IV  NOT_1392(II3923,n2710gat);
  IV  NOT_1393(n2707gat,II3923);
  IV  NOT_1394(n16gat,n564gat);
  IV  NOT_1395(n295gat,n357gat);
  IV  NOT_1396(n11gat,n12gat);
  IV  NOT_1397(n1889gat,n1961gat);
  IV  NOT_1398(II3935,n2704gat);
  IV  NOT_1399(n2700gat,II3935);
  IV  NOT_1400(n2051gat,n2056gat);
  IV  NOT_1401(II3941,n2684gat);
  IV  NOT_1402(n2680gat,II3941);
  IV  NOT_1403(n1350gat,n1831gat);
  IV  NOT_1404(II3945,n1350gat);
  IV  NOT_1405(n2696gat,II3945);
  IV  NOT_1406(II3948,n2696gat);
  IV  NOT_1407(n2692gat,II3948);
  IV  NOT_1408(II3951,n2448gat);
  IV  NOT_1409(n2683gat,II3951);
  IV  NOT_1410(II3954,n2683gat);
  IV  NOT_1411(n2679gat,II3954);
  IV  NOT_1412(II3957,n2450gat);
  IV  NOT_1413(n2449gat,II3957);
  IV  NOT_1414(n1754gat,n2449gat);
  IV  NOT_1415(II3962,n2830gat);
  IV  NOT_1416(n2827gat,II3962);
  IV  NOT_1417(n2590gat,n2592gat);
  IV  NOT_1418(n2456gat,n2458gat);
  IV  NOT_1419(n2512gat,n2514gat);
  IV  NOT_1420(n1544gat,n1625gat);
  IV  NOT_1421(n1769gat,n1771gat);
  IV  NOT_1422(n1683gat,n1756gat);
  IV  NOT_1423(n2167gat,n2169gat);
  IV  NOT_1424(n2013gat,II4000);
  IV  NOT_1425(n1791gat,n2013gat);
  IV  NOT_1426(n2691gat,n2695gat);
  IV  NOT_1427(n1518gat,n1694gat);
  IV  NOT_1428(n2699gat,n2703gat);
  IV  NOT_1429(n2159gat,n1412gat);
  IV  NOT_1430(n2478gat,n2579gat);
  IV  NOT_1431(II4014,n2744gat);
  IV  NOT_1432(n2740gat,II4014);
  IV  NOT_1433(n2158gat,n1412gat);
  IV  NOT_1434(n2186gat,n2613gat);
  IV  NOT_1435(II4020,n2800gat);
  IV  NOT_1436(n2797gat,II4020);
  IV  NOT_1437(n2288gat,II4024);
  IV  NOT_1438(n1513gat,n2288gat);
  IV  NOT_1439(n2537gat,n2538gat);
  IV  NOT_1440(n2442gat,n2483gat);
  IV  NOT_1441(n1334gat,n1336gat);
  IV  NOT_1442(II4055,n1748gat);
  IV  NOT_1443(n1747gat,II4055);
  IV  NOT_1444(II4067,n1675gat);
  IV  NOT_1445(n1674gat,II4067);
  IV  NOT_1446(n1403gat,n1402gat);
  IV  NOT_1447(II4081,n1807gat);
  IV  NOT_1448(n1806gat,II4081);
  IV  NOT_1449(n1634gat,n1712gat);
  IV  NOT_1450(n1338gat,n1340gat);
  IV  NOT_1451(II4105,n1456gat);
  IV  NOT_1452(n1455gat,II4105);
  IV  NOT_1453(II4108,n1340gat);
  IV  NOT_1454(n1339gat,II4108);
  IV  NOT_1455(n1505gat,n2980gat);
  IV  NOT_1456(II4117,n1505gat);
  IV  NOT_1457(n2758gat,II4117);
  IV  NOT_1458(n2755gat,n2758gat);
  IV  NOT_1459(n1546gat,n2980gat);
  IV  NOT_1460(II4122,n1546gat);
  IV  NOT_1461(n2752gat,II4122);
  IV  NOT_1462(n2748gat,n2752gat);
  IV  NOT_1463(n2012gat,n2016gat);
  IV  NOT_1464(n2002gat,n2008gat);
  IV  NOT_1465(II4129,n3097gat);
  IV  NOT_1466(n2858gat,II4129);
  IV  NOT_1467(n2857gat,n2858gat);
  IV  NOT_1468(II4135,n3098gat);
  IV  NOT_1469(n2766gat,II4135);
  IV  NOT_1470(II4138,n2766gat);
  IV  NOT_1471(n2765gat,II4138);
  IV  NOT_1472(n1684gat,n1759gat);
  IV  NOT_1473(n1632gat,II4145);
  IV  NOT_1474(II4157,n1525gat);
  IV  NOT_1475(n1524gat,II4157);
  IV  NOT_1476(n1862gat,n1863gat);
  IV  NOT_1477(n1919gat,n1860gat);
  IV  NOT_1478(n1460gat,n1462gat);
  IV  NOT_1479(II4185,n1596gat);
  IV  NOT_1480(n1595gat,II4185);
  IV  NOT_1481(n1454gat,n1469gat);
  IV  NOT_1482(n1468gat,n1519gat);
  IV  NOT_1483(II4194,n1462gat);
  IV  NOT_1484(n1461gat,II4194);
  IV  NOT_1485(n1477gat,n2984gat);
  IV  NOT_1486(n1594gat,n1596gat);
  IV  NOT_1487(II4212,n1588gat);
  IV  NOT_1488(n1587gat,II4212);
  IV  NOT_1489(n1681gat,II4217);
  IV  NOT_1490(II4222,n1761gat);
  IV  NOT_1491(n2751gat,II4222);
  IV  NOT_1492(n2747gat,n2751gat);
  IV  NOT_1493(II4227,n1760gat);
  IV  NOT_1494(n2743gat,II4227);
  IV  NOT_1495(n2739gat,n2743gat);
  IV  NOT_1496(n1978gat,n2286gat);
  IV  NOT_1497(II4233,n1721gat);
  IV  NOT_1498(n2808gat,II4233);
  IV  NOT_1499(II4236,n2808gat);
  IV  NOT_1500(n2804gat,II4236);
  IV  NOT_1501(n517gat,n518gat);
  IV  NOT_1502(n417gat,n418gat);
  IV  NOT_1503(n413gat,n411gat);
  IV  NOT_1504(n412gat,n522gat);
  IV  NOT_1505(n406gat,n516gat);
  IV  NOT_1506(n407gat,n355gat);
  IV  NOT_1507(n290gat,n525gat);
  IV  NOT_1508(n527gat,n356gat);
  IV  NOT_1509(n416gat,n415gat);
  IV  NOT_1510(n528gat,n521gat);
  IV  NOT_1511(n358gat,n532gat);
  IV  NOT_1512(n639gat,n523gat);
  IV  NOT_1513(n1111gat,n635gat);
  IV  NOT_1514(n524gat,n414gat);
  IV  NOT_1515(n1112gat,n630gat);
  IV  NOT_1516(n741gat,n629gat);
  IV  NOT_1517(n633gat,n634gat);
  IV  NOT_1518(n926gat,n632gat);
  IV  NOT_1519(n670gat,n636gat);
  IV  NOT_1520(n1123gat,n632gat);
  IV  NOT_1521(n1007gat,n635gat);
  IV  NOT_1522(n1006gat,n630gat);
  IV  NOT_1523(II4309,n2941gat);
  IV  NOT_1524(n2814gat,II4309);
  IV  NOT_1525(II4312,n2814gat);
  IV  NOT_1526(n2811gat,II4312);
  IV  NOT_1527(n1002gat,n2946gat);
  IV  NOT_1528(II4329,n2950gat);
  IV  NOT_1529(n2813gat,II4329);
  IV  NOT_1530(II4332,n2813gat);
  IV  NOT_1531(n2810gat,II4332);
  IV  NOT_1532(n888gat,n2933gat);
  IV  NOT_1533(II4349,n2935gat);
  IV  NOT_1534(n2818gat,II4349);
  IV  NOT_1535(II4352,n2818gat);
  IV  NOT_1536(n2816gat,II4352);
  IV  NOT_1537(n898gat,n2940gat);
  IV  NOT_1538(II4369,n2937gat);
  IV  NOT_1539(n2817gat,II4369);
  IV  NOT_1540(II4372,n2817gat);
  IV  NOT_1541(n2815gat,II4372);
  IV  NOT_1542(n1179gat,n2947gat);
  IV  NOT_1543(II4389,n2956gat);
  IV  NOT_1544(n2824gat,II4389);
  IV  NOT_1545(II4392,n2824gat);
  IV  NOT_1546(n2821gat,II4392);
  IV  NOT_1547(n897gat,n2939gat);
  IV  NOT_1548(II4409,n2938gat);
  IV  NOT_1549(n2823gat,II4409);
  IV  NOT_1550(II4412,n2823gat);
  IV  NOT_1551(n2820gat,II4412);
  IV  NOT_1552(n894gat,n2932gat);
  IV  NOT_1553(II4429,n2936gat);
  IV  NOT_1554(n2829gat,II4429);
  IV  NOT_1555(II4432,n2829gat);
  IV  NOT_1556(n2826gat,II4432);
  IV  NOT_1557(n1180gat,n2948gat);
  IV  NOT_1558(II4449,n2955gat);
  IV  NOT_1559(n2828gat,II4449);
  IV  NOT_1560(II4452,n2828gat);
  IV  NOT_1561(n2825gat,II4452);
  IV  NOT_1562(n671gat,n673gat);
  IV  NOT_1563(n628gat,n631gat);
  IV  NOT_1564(n976gat,n628gat);
  IV  NOT_1565(II4475,n2951gat);
  IV  NOT_1566(n2807gat,II4475);
  IV  NOT_1567(II4478,n2807gat);
  IV  NOT_1568(n2803gat,II4478);
  IV  NOT_1569(n2127gat,n2389gat);
  IV  NOT_1570(II4482,n2127gat);
  IV  NOT_1571(n2682gat,II4482);
  IV  NOT_1572(II4485,n2682gat);
  IV  NOT_1573(n2678gat,II4485);
  IV  NOT_1574(n2046gat,n2269gat);
  IV  NOT_1575(II4489,n2046gat);
  IV  NOT_1576(n2681gat,II4489);
  IV  NOT_1577(II4492,n2681gat);
  IV  NOT_1578(n2677gat,II4492);
  IV  NOT_1579(n1708gat,n2338gat);
  IV  NOT_1580(II4496,n1708gat);
  IV  NOT_1581(n2688gat,II4496);
  IV  NOT_1582(II4499,n2688gat);
  IV  NOT_1583(n2686gat,II4499);
  IV  NOT_1584(n455gat,n291gat);
  IV  NOT_1585(n2237gat,n2646gat);
  IV  NOT_1586(II4506,n2764gat);
  IV  NOT_1587(n2763gat,II4506);
  IV  NOT_1588(n1782gat,n2971gat);
  IV  NOT_1589(II4512,n2762gat);
  IV  NOT_1590(n2760gat,II4512);
  IV  NOT_1591(n2325gat,n3010gat);
  IV  NOT_1592(II4518,n2761gat);
  IV  NOT_1593(n2759gat,II4518);
  IV  NOT_1594(n2245gat,n504gat);
  IV  NOT_1595(II4524,n2757gat);
  IV  NOT_1596(n2754gat,II4524);
  IV  NOT_1597(n2244gat,n567gat);
  IV  NOT_1598(II4530,n2756gat);
  IV  NOT_1599(n2753gat,II4530);
  IV  NOT_1600(n2243gat,n55gat);
  IV  NOT_1601(II4536,n2750gat);
  IV  NOT_1602(n2746gat,II4536);
  IV  NOT_1603(n2246gat,n933gat);
  IV  NOT_1604(II4542,n2749gat);
  IV  NOT_1605(n2745gat,II4542);
  IV  NOT_1606(n2384gat,n43gat);
  IV  NOT_1607(II4548,n2742gat);
  IV  NOT_1608(n2738gat,II4548);
  IV  NOT_1609(n2385gat,n748gat);
  IV  NOT_1610(II4554,n2741gat);
  IV  NOT_1611(n2737gat,II4554);
  IV  NOT_1612(n1286gat,n1269gat);
  IV  NOT_1613(II4558,n1286gat);
  IV  NOT_1614(n2687gat,II4558);
  IV  NOT_1615(n2685gat,n2687gat);
  IV  NOT_1616(n1328gat,n1224gat);
  IV  NOT_1617(n1381gat,n1328gat);
  IV  NOT_1618(n1384gat,n2184gat);
  IV  NOT_1619(II4566,n2694gat);
  IV  NOT_1620(n2690gat,II4566);
  IV  NOT_1621(n1382gat,n1280gat);
  IV  NOT_1622(n1451gat,n1382gat);
  IV  NOT_1623(n1453gat,n2187gat);
  IV  NOT_1624(II4573,n2693gat);
  IV  NOT_1625(n2689gat,II4573);
  IV  NOT_1626(n927gat,n1133gat);
  IV  NOT_1627(n925gat,n927gat);
  IV  NOT_1628(n1452gat,n2049gat);
  IV  NOT_1629(II4580,n2702gat);
  IV  NOT_1630(n2698gat,II4580);
  IV  NOT_1631(n923gat,n1043gat);
  IV  NOT_1632(n921gat,n923gat);
  IV  NOT_1633(n1890gat,n2328gat);
  IV  NOT_1634(II4587,n2701gat);
  IV  NOT_1635(n2697gat,II4587);
  IV  NOT_1636(n850gat,n929gat);
  IV  NOT_1637(n739gat,n850gat);
  IV  NOT_1638(n1841gat,n2058gat);
  IV  NOT_1639(II4594,n2709gat);
  IV  NOT_1640(n2706gat,II4594);
  IV  NOT_1641(n922gat,n1119gat);
  IV  NOT_1642(n848gat,n922gat);
  IV  NOT_1643(n2047gat,n2209gat);
  IV  NOT_1644(II4601,n2708gat);
  IV  NOT_1645(n2705gat,II4601);
  IV  NOT_1646(n924gat,n1070gat);
  IV  NOT_1647(n849gat,n924gat);
  IV  NOT_1648(n2050gat,n2146gat);
  IV  NOT_1649(II4608,n2799gat);
  IV  NOT_1650(n2796gat,II4608);
  IV  NOT_1651(n1118gat,n1033gat);
  IV  NOT_1652(n1032gat,n1118gat);
  IV  NOT_1653(n2054gat,n2281gat);
  IV  NOT_1654(II4615,n2798gat);
  IV  NOT_1655(n2795gat,II4615);
  IV  NOT_1656(II4620,n1745gat);
  IV  NOT_1657(n2806gat,II4620);
  IV  NOT_1658(II4623,n2806gat);
  IV  NOT_1659(n2802gat,II4623);
  IV  NOT_1660(II4626,n1871gat);
  IV  NOT_1661(n1870gat,II4626);
  IV  NOT_1662(n1086gat,n1870gat);
  IV  NOT_1663(II4630,n1086gat);
  IV  NOT_1664(n2805gat,II4630);
  IV  NOT_1665(II4633,n2805gat);
  IV  NOT_1666(n2801gat,II4633);
  IV  NOT_1667(n67gat,n85gat);
  IV  NOT_1668(n71gat,n180gat);
  IV  NOT_1669(n1840gat,n1892gat);
  IV  NOT_1670(II4642,n2812gat);
  IV  NOT_1671(n2809gat,II4642);
  IV  NOT_1672(n76gat,n82gat);
  IV  NOT_1673(n14gat,n186gat);
  IV  NOT_1674(n1842gat,n1711gat);
  IV  NOT_1675(II4651,n2822gat);
  IV  NOT_1676(n2819gat,II4651);
  IV  NOT_1677(II4654,n2819gat);
  IV  NOT_1678(n3104gat,II4654);
  IV  NOT_1679(II4657,n2809gat);
  IV  NOT_1680(n3105gat,II4657);
  IV  NOT_1681(II4660,n2801gat);
  IV  NOT_1682(n3106gat,II4660);
  IV  NOT_1683(II4663,n2802gat);
  IV  NOT_1684(n3107gat,II4663);
  IV  NOT_1685(II4666,n2795gat);
  IV  NOT_1686(n3108gat,II4666);
  IV  NOT_1687(II4669,n2796gat);
  IV  NOT_1688(n3109gat,II4669);
  IV  NOT_1689(II4672,n2705gat);
  IV  NOT_1690(n3110gat,II4672);
  IV  NOT_1691(II4675,n2706gat);
  IV  NOT_1692(n3111gat,II4675);
  IV  NOT_1693(II4678,n2697gat);
  IV  NOT_1694(n3112gat,II4678);
  IV  NOT_1695(II4681,n2698gat);
  IV  NOT_1696(n3113gat,II4681);
  IV  NOT_1697(II4684,n2689gat);
  IV  NOT_1698(n3114gat,II4684);
  IV  NOT_1699(II4687,n2690gat);
  IV  NOT_1700(n3115gat,II4687);
  IV  NOT_1701(II4690,n2685gat);
  IV  NOT_1702(n3116gat,II4690);
  IV  NOT_1703(II4693,n2737gat);
  IV  NOT_1704(n3117gat,II4693);
  IV  NOT_1705(II4696,n2738gat);
  IV  NOT_1706(n3118gat,II4696);
  IV  NOT_1707(II4699,n2745gat);
  IV  NOT_1708(n3119gat,II4699);
  IV  NOT_1709(II4702,n2746gat);
  IV  NOT_1710(n3120gat,II4702);
  IV  NOT_1711(II4705,n2753gat);
  IV  NOT_1712(n3121gat,II4705);
  IV  NOT_1713(II4708,n2754gat);
  IV  NOT_1714(n3122gat,II4708);
  IV  NOT_1715(II4711,n2759gat);
  IV  NOT_1716(n3123gat,II4711);
  IV  NOT_1717(II4714,n2760gat);
  IV  NOT_1718(n3124gat,II4714);
  IV  NOT_1719(II4717,n2763gat);
  IV  NOT_1720(n3125gat,II4717);
  IV  NOT_1721(II4720,n2686gat);
  IV  NOT_1722(n3126gat,II4720);
  IV  NOT_1723(II4723,n2677gat);
  IV  NOT_1724(n3127gat,II4723);
  IV  NOT_1725(II4726,n2678gat);
  IV  NOT_1726(n3128gat,II4726);
  IV  NOT_1727(II4729,n2803gat);
  IV  NOT_1728(n3129gat,II4729);
  IV  NOT_1729(II4732,n2825gat);
  IV  NOT_1730(n3130gat,II4732);
  IV  NOT_1731(II4735,n2826gat);
  IV  NOT_1732(n3131gat,II4735);
  IV  NOT_1733(II4738,n2820gat);
  IV  NOT_1734(n3132gat,II4738);
  IV  NOT_1735(II4741,n2821gat);
  IV  NOT_1736(n3133gat,II4741);
  IV  NOT_1737(II4744,n2815gat);
  IV  NOT_1738(n3134gat,II4744);
  IV  NOT_1739(II4747,n2816gat);
  IV  NOT_1740(n3135gat,II4747);
  IV  NOT_1741(II4750,n2810gat);
  IV  NOT_1742(n3136gat,II4750);
  IV  NOT_1743(II4753,n2811gat);
  IV  NOT_1744(n3137gat,II4753);
  IV  NOT_1745(II4756,n2804gat);
  IV  NOT_1746(n3138gat,II4756);
  IV  NOT_1747(II4759,n2739gat);
  IV  NOT_1748(n3139gat,II4759);
  IV  NOT_1749(II4762,n2747gat);
  IV  NOT_1750(n3140gat,II4762);
  IV  NOT_1751(II4765,n2748gat);
  IV  NOT_1752(n3141gat,II4765);
  IV  NOT_1753(II4768,n2755gat);
  IV  NOT_1754(n3142gat,II4768);
  IV  NOT_1755(II4771,n2797gat);
  IV  NOT_1756(n3143gat,II4771);
  IV  NOT_1757(II4774,n2740gat);
  IV  NOT_1758(n3144gat,II4774);
  IV  NOT_1759(II4777,n2699gat);
  IV  NOT_1760(n3145gat,II4777);
  IV  NOT_1761(II4780,n2691gat);
  IV  NOT_1762(n3146gat,II4780);
  IV  NOT_1763(II4783,n2827gat);
  IV  NOT_1764(n3147gat,II4783);
  IV  NOT_1765(II4786,n2679gat);
  IV  NOT_1766(n3148gat,II4786);
  IV  NOT_1767(II4789,n2692gat);
  IV  NOT_1768(n3149gat,II4789);
  IV  NOT_1769(II4792,n2680gat);
  IV  NOT_1770(n3150gat,II4792);
  IV  NOT_1771(II4795,n2700gat);
  IV  NOT_1772(n3151gat,II4795);
  IV  NOT_1773(II4798,n2707gat);
  IV  NOT_1774(n3152gat,II4798);
  OR2 OR2_0(n2897gat,n648gat,n442gat);
  OR4 OR4_0(n1213gat,n1214gat,n1215gat,n1216gat,n1217gat);
  OR2 OR2_1(n2906gat,n745gat,n638gat);
  OR2 OR2_2(n2889gat,n423gat,n362gat);
  OR4 OR4_1(n748gat,n749gat,n750gat,n751gat,n752gat);
  OR4 OR4_2(n258gat,n259gat,n260gat,n261gat,n262gat);
  OR4 OR4_3(n1013gat,n1014gat,n1015gat,n1016gat,n1017gat);
  OR4 OR4_4(n475gat,n476gat,n477gat,n478gat,n479gat);
  OR4 OR4_5(n43gat,n44gat,n45gat,n46gat,n47gat);
  OR2 OR2_3(n2786gat,n3091gat,n3092gat);
  OR4 OR4_6(n167gat,n168gat,n169gat,n170gat,n171gat);
  OR4 OR4_7(n906gat,n907gat,n908gat,n909gat,n910gat);
  OR4 OR4_8(n343gat,n344gat,n345gat,n346gat,n347gat);
  OR4 OR4_9(n55gat,n56gat,n57gat,n58gat,n59gat);
  OR2 OR2_4(n2914gat,n768gat,n655gat);
  OR2 OR2_5(n2928gat,n963gat,n868gat);
  OR2 OR2_6(n2927gat,n962gat,n959gat);
  OR4 OR4_10(n944gat,n945gat,n946gat,n947gat,n948gat);
  OR2 OR2_7(n2896gat,n647gat,n441gat);
  OR2 OR2_8(n2922gat,n967gat,n792gat);
  OR4 OR4_11(n1228gat,n1229gat,n1230gat,n1231gat,n1232gat);
  OR2 OR2_9(n2894gat,n443gat,n439gat);
  OR2 OR2_10(n2921gat,n966gat,n790gat);
  OR2 OR2_11(n2895gat,n444gat,n440gat);
  OR4 OR4_12(n1050gat,n1051gat,n1052gat,n1053gat,n1054gat);
  OR4 OR4_13(n933gat,n934gat,n935gat,n936gat,n937gat);
  OR4 OR4_14(n709gat,n710gat,n711gat,n712gat,n713gat);
  OR4 OR4_15(n728gat,n729gat,n730gat,n731gat,n732gat);
  OR4 OR4_16(n493gat,n494gat,n495gat,n496gat,n497gat);
  OR4 OR4_17(n504gat,n505gat,n506gat,n507gat,n508gat);
  OR3 OR3_0(II1277,n2860gat,n2855gat,n2863gat);
  OR3 OR3_1(II1278,n740gat,n3030gat,II1277);
  OR2 OR2_12(n2913gat,n767gat,n653gat);
  OR2 OR2_13(n2920gat,n867gat,n771gat);
  OR2 OR2_14(n2905gat,n964gat,n961gat);
  OR4 OR4_18(n803gat,n804gat,n805gat,n806gat,n807gat);
  OR4 OR4_19(n586gat,n587gat,n588gat,n589gat,n590gat);
  OR2 OR2_15(n2898gat,n447gat,n445gat);
  OR4 OR4_20(n686gat,n687gat,n688gat,n689gat,n690gat);
  OR4 OR4_21(n567gat,n568gat,n569gat,n570gat,n571gat);
  OR3 OR3_2(II1515,n2474gat,n2524gat,n2831gat);
  OR3 OR3_3(II1516,n2466gat,n2462gat,II1515);
  OR3 OR3_4(II1584,n2353gat,n2284gat,n2354gat);
  OR3 OR3_5(II1585,n2356gat,n2214gat,II1584);
  OR2 OR2_16(n2989gat,n1693gat,n1692gat);
  OR3 OR3_6(II1723,n2354gat,n2353gat,n2214gat);
  OR3 OR3_7(II1724,n2355gat,n2443gat,II1723);
  OR3 OR3_8(II1733,n2286gat,n2428gat,n2289gat);
  OR3 OR3_9(II1734,n1604gat,n2214gat,II1733);
  OR2 OR2_17(n2918gat,n769gat,n759gat);
  OR2 OR2_18(n2952gat,n1076gat,n1075gat);
  OR2 OR2_19(n2919gat,n766gat,n760gat);
  OR4 OR4_22(n1184gat,n1185gat,n1186gat,n1187gat,n1188gat);
  OR2 OR2_20(n2910gat,n645gat,n644gat);
  OR2 OR2_21(n2907gat,n646gat,n641gat);
  OR2 OR2_22(n2970gat,n1383gat,n1327gat);
  OR2 OR2_23(n2911gat,n761gat,n651gat);
  OR2 OR2_24(n2912gat,n762gat,n652gat);
  OR2 OR2_25(n2909gat,n765gat,n643gat);
  OR4 OR4_23(n1201gat,n1202gat,n1203gat,n1204gat,n1205gat);
  OR4 OR4_24(n1269gat,n1270gat,n1271gat,n1272gat,n1273gat);
  OR2 OR2_26(n2908gat,n763gat,n642gat);
  OR2 OR2_27(n2971gat,n1287gat,n1285gat);
  OR3 OR3_10(n2904gat,n793gat,n664gat,n556gat);
  OR3 OR3_11(n2891gat,n795gat,n656gat,n368gat);
  OR3 OR3_12(n2903gat,n794gat,n773gat,n662gat);
  OR3 OR3_13(n2915gat,n965gat,n960gat,n661gat);
  OR4 OR4_25(n779gat,n780gat,n781gat,n782gat,n783gat);
  OR3 OR3_14(n2901gat,n558gat,n555gat,n450gat);
  OR3 OR3_15(n2890gat,n654gat,n557gat,n371gat);
  OR2 OR2_28(n2876gat,n874gat,n132gat);
  OR3 OR3_16(n2888gat,n663gat,n649gat,n449gat);
  OR3 OR3_17(n2887gat,n791gat,n650gat,n370gat);
  OR3 OR3_18(n2886gat,n774gat,n764gat,n369gat);
  OR4 OR4_26(n221gat,n222gat,n223gat,n224gat,n225gat);
  OR4 OR4_27(n120gat,n121gat,n122gat,n123gat,n124gat);
  OR2 OR2_29(n3010gat,n2460gat,n2423gat);
  OR2 OR2_30(n3016gat,n2596gat,n2595gat);
  OR4 OR4_28(n2568gat,n2569gat,n2570gat,n2571gat,n2572gat);
  OR4 OR4_29(n2409gat,n2410gat,n2411gat,n2412gat,n2413gat);
  OR2 OR2_31(n2579gat,n2580gat,n2581gat);
  OR2 OR2_32(n3014gat,n2567gat,n2499gat);
  OR2 OR2_33(n2880gat,n299gat,n207gat);
  OR2 OR2_34(n2646gat,n2647gat,n2648gat);
  OR4 OR4_30(n2601gat,n2602gat,n2603gat,n2604gat,n2605gat);
  OR4 OR4_31(n2545gat,n2546gat,n2547gat,n2548gat,n2549gat);
  OR2 OR2_35(n2613gat,n2614gat,n2615gat);
  OR2 OR2_36(n3013gat,n2461gat,n2421gat);
  OR4 OR4_32(n2930gat,n1153gat,n1151gat,n982gat,n877gat);
  OR4 OR4_33(n2957gat,n1159gat,n1158gat,n1156gat,n1155gat);
  OR2 OR2_37(n2975gat,n1443gat,n1325gat);
  OR2 OR2_38(n2974gat,n1321gat,n1320gat);
  OR2 OR2_39(n2966gat,n1368gat,n1258gat);
  OR2 OR2_40(n2979gat,n1373gat,n1372gat);
  OR4 OR4_34(n2978gat,n1441gat,n1440gat,n1371gat,n1367gat);
  OR2 OR2_41(n2982gat,n1504gat,n1502gat);
  OR2 OR2_42(n2954gat,n1250gat,n1103gat);
  OR2 OR2_43(n2964gat,n1304gat,n1249gat);
  OR2 OR2_44(n2958gat,n1246gat,n1161gat);
  OR2 OR2_45(n2963gat,n1291gat,n1245gat);
  OR4 OR4_35(n2973gat,n1352gat,n1351gat,n1303gat,n1302gat);
  OR2 OR2_46(n2953gat,n1163gat,n1102gat);
  OR2 OR2_47(n2949gat,n1101gat,n996gat);
  OR2 OR2_48(n2934gat,n1104gat,n887gat);
  OR2 OR2_49(n2959gat,n1305gat,n1162gat);
  OR4 OR4_36(n2977gat,n1360gat,n1359gat,n1358gat,n1357gat);
  OR3 OR3_19(II2720,n1788gat,n1786gat,n1839gat);
  OR3 OR3_20(II2721,n1884gat,n1783gat,II2720);
  OR3 OR3_21(II2735,n1788gat,n1884gat,n1633gat);
  OR3 OR3_22(II2736,n1785gat,n1784gat,II2735);
  OR3 OR3_23(II2812,n1703gat,n1704gat,n1778gat);
  OR4 OR4_37(II2813,n1609gat,n1702gat,n1700gat,II2812);
  OR3 OR3_24(II2831,n1839gat,n1786gat,n1788gat);
  OR3 OR3_25(II2832,n1884gat,n1784gat,II2831);
  OR3 OR3_26(II2889,n1784gat,n1633gat,n1884gat);
  OR3 OR3_27(II2890,n1788gat,n1786gat,II2889);
  OR3 OR3_28(II2925,n1784gat,n1785gat,n1633gat);
  OR3 OR3_29(II2926,n1884gat,n1787gat,II2925);
  OR3 OR3_30(II2934,n1784gat,n1839gat,n1788gat);
  OR3 OR3_31(II2935,n1785gat,n1884gat,II2934);
  OR2 OR2_50(n2988gat,n1733gat,n1581gat);
  OR2 OR2_51(n2983gat,n2079gat,n2073gat);
  OR2 OR2_52(n2987gat,n1574gat,n1573gat);
  OR3 OR3_32(n2992gat,n1723gat,n1647gat,n1646gat);
  OR3 OR3_33(n2986gat,n1650gat,n1649gat,n1563gat);
  OR3 OR3_34(n2991gat,n1654gat,n1653gat,n1644gat);
  OR3 OR3_35(II3148,n1839gat,n1884gat,n1784gat);
  OR3 OR3_36(II3149,n1786gat,n1787gat,II3148);
  OR3 OR3_37(II3178,n1838gat,n1785gat,n1788gat);
  OR3 OR3_38(II3179,n1839gat,n1784gat,II3178);
  OR3 OR3_39(n2981gat,n1413gat,n1408gat,n1407gat);
  OR2 OR2_53(n3000gat,n2000gat,n1999gat);
  OR3 OR3_40(n3004gat,n2258gat,n2257gat,n2255gat);
  OR2 OR2_54(n3003gat,n2256gat,n2251gat);
  OR2 OR2_55(n3001gat,n2132gat,n2130gat);
  OR2 OR2_56(n3006gat,n2253gat,n2252gat);
  OR2 OR2_57(n3007gat,n2250gat,n2249gat);
  OR2 OR2_58(n2990gat,n1710gat,n1630gat);
  OR2 OR2_59(n2994gat,n1954gat,n1888gat);
  OR3 OR3_41(n2993gat,n1894gat,n1847gat,n1846gat);
  OR2 OR2_60(n2998gat,n2055gat,n1967gat);
  OR3 OR3_42(n2996gat,n1960gat,n1959gat,n1957gat);
  OR2 OR2_61(n3008gat,n2332gat,n2259gat);
  OR2 OR2_62(n3005gat,n2211gat,n2210gat);
  OR3 OR3_43(n2997gat,n2053gat,n2052gat,n1964gat);
  OR2 OR2_63(n3009gat,n2350gat,n2282gat);
  OR3 OR3_44(n3002gat,n2213gat,n2150gat,n2149gat);
  OR2 OR2_64(n2995gat,n1962gat,n1955gat);
  OR2 OR2_65(n2999gat,n1972gat,n1971gat);
  OR2 OR2_66(n3011gat,n2333gat,n2331gat);
  OR2 OR2_67(n3015gat,n2566gat,n2565gat);
  OR3 OR3_45(n2874gat,n141gat,n38gat,n37gat);
  OR2 OR2_68(n2917gat,n1074gat,n872gat);
  OR2 OR2_69(n2878gat,n234gat,n137gat);
  OR2 OR2_70(n2892gat,n378gat,n377gat);
  OR3 OR3_46(n2885gat,n250gat,n249gat,n248gat);
  OR3 OR3_47(n2900gat,n869gat,n453gat,n448gat);
  OR2 OR2_71(n2883gat,n251gat,n244gat);
  OR3 OR3_48(n2929gat,n974gat,n973gat,n870gat);
  OR2 OR2_72(n2884gat,n246gat,n245gat);
  OR2 OR2_73(n2902gat,n460gat,n459gat);
  OR3 OR3_49(n2925gat,n975gat,n972gat,n969gat);
  OR2 OR2_74(n2879gat,n145gat,n143gat);
  OR3 OR3_50(n2916gat,n971gat,n970gat,n968gat);
  OR3 OR3_51(n2875gat,n142gat,n40gat,n39gat);
  OR3 OR3_52(n2899gat,n772gat,n451gat,n446gat);
  OR2 OR2_75(n2877gat,n139gat,n136gat);
  OR2 OR2_76(n2893gat,n391gat,n390gat);
  OR2 OR2_77(n2926gat,n1083gat,n1077gat);
  OR2 OR2_78(n2882gat,n242gat,n240gat);
  OR2 OR2_79(n2924gat,n871gat,n797gat);
  OR3 OR3_53(n2881gat,n324gat,n238gat,n237gat);
  OR2 OR2_80(n2923gat,n1082gat,n796gat);
  OR2 OR2_81(n2710gat,n69gat,n1885gat);
  OR2 OR2_82(n2704gat,n11gat,n1889gat);
  OR2 OR2_83(n2684gat,n1599gat,n2051gat);
  OR2 OR2_84(n2830gat,n2444gat,n1754gat);
  OR3 OR3_54(II3999,n2167gat,n2031gat,n2174gat);
  OR4 OR4_38(II4000,n2108gat,n2093gat,n2035gat,II3999);
  OR2 OR2_85(n2695gat,n1586gat,n1791gat);
  OR2 OR2_86(n2703gat,n1755gat,n1518gat);
  OR2 OR2_87(n2744gat,n2159gat,n2478gat);
  OR2 OR2_88(n2800gat,n2158gat,n2186gat);
  OR3 OR3_55(II4023,n2443gat,n2290gat,n2214gat);
  OR3 OR3_56(II4024,n2353gat,n2284gat,II4023);
  OR4 OR4_39(n2980gat,n1470gat,n1400gat,n1399gat,n1398gat);
  OR3 OR3_57(II4144,n1633gat,n1838gat,n1786gat);
  OR3 OR3_58(II4145,n1788gat,n1784gat,II4144);
  OR2 OR2_89(n2984gat,n1467gat,n1466gat);
  OR4 OR4_40(n2985gat,n1686gat,n1533gat,n1532gat,n1531gat);
  OR3 OR3_59(II4216,n1427gat,n1595gat,n1677gat);
  OR3 OR3_60(II4217,n1392gat,n2989gat,II4216);
  OR4 OR4_41(n2931gat,n1100gat,n994gat,n989gat,n880gat);
  OR2 OR2_90(n2943gat,n1012gat,n905gat);
  OR2 OR2_91(n2941gat,n1003gat,n902gat);
  OR4 OR4_42(n2946gat,n1099gat,n998gat,n995gat,n980gat);
  OR2 OR2_92(n2960gat,n1175gat,n1174gat);
  OR2 OR2_93(n2950gat,n1001gat,n999gat);
  OR2 OR2_94(n2969gat,n1323gat,n1264gat);
  OR4 OR4_43(n2933gat,n981gat,n890gat,n889gat,n886gat);
  OR2 OR2_95(n2935gat,n892gat,n891gat);
  OR2 OR2_96(n2942gat,n904gat,n903gat);
  OR4 OR4_44(n2940gat,n1152gat,n1092gat,n997gat,n993gat);
  OR2 OR2_97(n2937gat,n900gat,n895gat);
  OR4 OR4_45(n2947gat,n1094gat,n1093gat,n988gat,n984gat);
  OR2 OR2_98(n2965gat,n1267gat,n1257gat);
  OR2 OR2_99(n2956gat,n1178gat,n1116gat);
  OR2 OR2_100(n2961gat,n1375gat,n1324gat);
  OR4 OR4_46(n2939gat,n1091gat,n1088gat,n992gat,n987gat);
  OR2 OR2_101(n2938gat,n899gat,n896gat);
  OR2 OR2_102(n2967gat,n1262gat,n1260gat);
  OR4 OR4_47(n2932gat,n1098gat,n1090gat,n986gat,n885gat);
  OR2 OR2_103(n2936gat,n901gat,n893gat);
  OR4 OR4_48(n2948gat,n1097gat,n1089gat,n1087gat,n991gat);
  OR2 OR2_104(n2968gat,n1326gat,n1261gat);
  OR2 OR2_105(n2955gat,n1177gat,n1115gat);
  OR2 OR2_106(n2944gat,n977gat,n976gat);
  OR4 OR4_49(n2945gat,n1096gat,n1095gat,n990gat,n979gat);
  OR2 OR2_107(n2962gat,n1176gat,n1173gat);
  OR2 OR2_108(n2951gat,n1004gat,n1000gat);
  OR2 OR2_109(n2764gat,n1029gat,n2237gat);
  OR2 OR2_110(n2762gat,n1028gat,n1782gat);
  OR2 OR2_111(n2761gat,n1031gat,n2325gat);
  OR2 OR2_112(n2757gat,n1030gat,n2245gat);
  OR2 OR2_113(n2756gat,n1011gat,n2244gat);
  OR2 OR2_114(n2750gat,n1181gat,n2243gat);
  OR2 OR2_115(n2749gat,n1010gat,n2246gat);
  OR2 OR2_116(n2742gat,n1005gat,n2384gat);
  OR2 OR2_117(n2741gat,n1182gat,n2385gat);
  OR2 OR2_118(n2694gat,n1381gat,n1384gat);
  OR2 OR2_119(n2693gat,n1451gat,n1453gat);
  OR2 OR2_120(n2702gat,n925gat,n1452gat);
  OR2 OR2_121(n2701gat,n921gat,n1890gat);
  OR2 OR2_122(n2709gat,n739gat,n1841gat);
  OR2 OR2_123(n2708gat,n848gat,n2047gat);
  OR2 OR2_124(n2799gat,n849gat,n2050gat);
  OR2 OR2_125(n2798gat,n1032gat,n2054gat);
  OR3 OR3_61(n2812gat,n73gat,n70gat,n1840gat);
  OR3 OR3_62(n2822gat,n77gat,n13gat,n1842gat);
  NR2 NOR2_0(n421gat,n2715gat,n2723gat);
  NR2 NOR2_1(n648gat,n373gat,n2669gat);
  NR2 NOR2_2(n442gat,n2844gat,n856gat);
  NR2 NOR2_3(n1499gat,n396gat,n401gat);
  NR2 NOR2_4(n1616gat,n918gat,n396gat);
  NR2 NOR2_5(n1614gat,n396gat,n845gat);
  NR3 NOR3_0(n1641gat,n1645gat,n1553gat,n1559gat);
  NR3 NOR3_1(n1642gat,n1559gat,n1616gat,n1645gat);
  NR3 NOR3_2(n1556gat,n1614gat,n1645gat,n1616gat);
  NR3 NOR3_3(n1557gat,n1553gat,n1645gat,n1614gat);
  NR3 NOR3_4(n1639gat,n1499gat,n1559gat,n1553gat);
  NR4 NOR4_0(n1605gat,n1614gat,n1616gat,n1499gat,n396gat);
  NR3 NOR3_5(n1555gat,n1616gat,n1559gat,n1499gat);
  NR3 NOR3_6(n1558gat,n1614gat,n1553gat,n1499gat);
  NR2 NOR2_6(n1256gat,n392gat,n702gat);
  NR2 NOR2_7(n1117gat,n720gat,n725gat);
  NR2 NOR2_8(n1618gat,n1319gat,n1447gat);
  NR2 NOR2_9(n1114gat,n725gat,n721gat);
  NR2 NOR2_10(n1621gat,n1319gat,n1380gat);
  NR2 NOR2_11(n1318gat,n392gat,n701gat);
  NR2 NOR2_12(n1619gat,n1447gat,n1446gat);
  NR2 NOR2_13(n1622gat,n1380gat,n1446gat);
  NR3 NOR3_7(n1214gat,n1218gat,n1219gat,n1220gat);
  NR3 NOR3_8(n1215gat,n1218gat,n1221gat,n1222gat);
  NR3 NOR3_9(n1216gat,n1223gat,n1219gat,n1222gat);
  NR3 NOR3_10(n1217gat,n1223gat,n1221gat,n1220gat);
  NR2 NOR2_14(n745gat,n2716gat,n2867gat);
  NR2 NOR2_15(n638gat,n2715gat,n2868gat);
  NR2 NOR2_16(n423gat,n2724gat,n2726gat);
  NR2 NOR2_17(n362gat,n2723gat,n2727gat);
  NR3 NOR3_11(n749gat,n753gat,n754gat,n755gat);
  NR3 NOR3_12(n750gat,n753gat,n756gat,n757gat);
  NR3 NOR3_13(n751gat,n758gat,n754gat,n757gat);
  NR3 NOR3_14(n752gat,n758gat,n756gat,n755gat);
  NR3 NOR3_15(n259gat,n263gat,n264gat,n265gat);
  NR3 NOR3_16(n260gat,n263gat,n266gat,n267gat);
  NR3 NOR3_17(n261gat,n268gat,n264gat,n267gat);
  NR3 NOR3_18(n262gat,n268gat,n266gat,n265gat);
  NR3 NOR3_19(n1014gat,n1018gat,n1019gat,n1020gat);
  NR3 NOR3_20(n1015gat,n1018gat,n1021gat,n1022gat);
  NR3 NOR3_21(n1016gat,n1023gat,n1019gat,n1022gat);
  NR3 NOR3_22(n1017gat,n1023gat,n1021gat,n1020gat);
  NR3 NOR3_23(n476gat,n480gat,n481gat,n482gat);
  NR3 NOR3_24(n477gat,n480gat,n483gat,n484gat);
  NR3 NOR3_25(n478gat,n485gat,n481gat,n484gat);
  NR3 NOR3_26(n479gat,n485gat,n483gat,n482gat);
  NR3 NOR3_27(n44gat,n48gat,n49gat,n50gat);
  NR3 NOR3_28(n45gat,n48gat,n51gat,n52gat);
  NR3 NOR3_29(n46gat,n53gat,n49gat,n52gat);
  NR3 NOR3_30(n47gat,n53gat,n51gat,n50gat);
  NR2 NOR2_18(n1376gat,n724gat,n720gat);
  NR2 NOR2_19(n1617gat,n1319gat,n1448gat);
  NR2 NOR2_20(n1377gat,n724gat,n721gat);
  NR2 NOR2_21(n1624gat,n1319gat,n1379gat);
  NR2 NOR2_22(n1113gat,n393gat,n701gat);
  NR2 NOR2_23(n1501gat,n1448gat,n1500gat);
  NR2 NOR2_24(n1623gat,n1379gat,n1446gat);
  NR2 NOR2_25(n1620gat,n1448gat,n1446gat);
  NR2 NOR2_26(n1827gat,n2729gat,n2317gat);
  NR2 NOR2_27(n1817gat,n1819gat,n1823gat);
  NR2 NOR2_28(n1935gat,n1816gat,n1828gat);
  NR2 NOR2_29(n529gat,n2724gat,n2715gat);
  NR2 NOR2_30(n361gat,n2859gat,n2726gat);
  NR3 NOR3_31(n168gat,n172gat,n173gat,n174gat);
  NR3 NOR3_32(n169gat,n172gat,n175gat,n176gat);
  NR3 NOR3_33(n170gat,n177gat,n173gat,n176gat);
  NR3 NOR3_34(n171gat,n177gat,n175gat,n174gat);
  NR3 NOR3_35(n907gat,n911gat,n912gat,n913gat);
  NR3 NOR3_36(n908gat,n911gat,n914gat,n915gat);
  NR3 NOR3_37(n909gat,n916gat,n912gat,n915gat);
  NR3 NOR3_38(n910gat,n916gat,n914gat,n913gat);
  NR3 NOR3_39(n344gat,n348gat,n349gat,n350gat);
  NR3 NOR3_40(n345gat,n348gat,n351gat,n352gat);
  NR3 NOR3_41(n346gat,n353gat,n349gat,n352gat);
  NR3 NOR3_42(n347gat,n353gat,n351gat,n350gat);
  NR3 NOR3_43(n56gat,n60gat,n61gat,n62gat);
  NR3 NOR3_44(n57gat,n60gat,n63gat,n64gat);
  NR3 NOR3_45(n58gat,n65gat,n61gat,n64gat);
  NR3 NOR3_46(n59gat,n65gat,n63gat,n62gat);
  NR2 NOR2_31(n768gat,n373gat,n2731gat);
  NR2 NOR2_32(n655gat,n856gat,n2718gat);
  NR2 NOR2_33(n963gat,n856gat,n2838gat);
  NR2 NOR2_34(n868gat,n2775gat,n373gat);
  NR2 NOR2_35(n962gat,n856gat,n2711gat);
  NR2 NOR2_36(n959gat,n373gat,n2734gat);
  NR3 NOR3_47(n945gat,n949gat,n950gat,n951gat);
  NR3 NOR3_48(n946gat,n949gat,n952gat,n953gat);
  NR3 NOR3_49(n947gat,n954gat,n950gat,n953gat);
  NR3 NOR3_50(n948gat,n954gat,n952gat,n951gat);
  NR2 NOR2_37(n647gat,n2792gat,n373gat);
  NR2 NOR2_38(n441gat,n856gat,n2846gat);
  NR2 NOR2_39(n967gat,n373gat,n2672gat);
  NR2 NOR2_40(n792gat,n2852gat,n856gat);
  NR3 NOR3_51(n1229gat,n1233gat,n1234gat,n1235gat);
  NR3 NOR3_52(n1230gat,n1233gat,n1236gat,n1237gat);
  NR3 NOR3_53(n1231gat,n1238gat,n1234gat,n1237gat);
  NR3 NOR3_54(n1232gat,n1238gat,n1236gat,n1235gat);
  NR2 NOR2_41(n443gat,n2778gat,n373gat);
  NR2 NOR2_42(n439gat,n856gat,n2836gat);
  NR2 NOR2_43(n966gat,n2789gat,n373gat);
  NR2 NOR2_44(n790gat,n856gat,n2840gat);
  NR2 NOR2_45(n444gat,n373gat,n2781gat);
  NR2 NOR2_46(n440gat,n856gat,n2842gat);
  NR3 NOR3_55(n1051gat,n1055gat,n1056gat,n1057gat);
  NR3 NOR3_56(n1052gat,n1055gat,n1058gat,n1059gat);
  NR3 NOR3_57(n1053gat,n1060gat,n1056gat,n1059gat);
  NR3 NOR3_58(n1054gat,n1060gat,n1058gat,n1057gat);
  NR3 NOR3_59(n934gat,n938gat,n939gat,n940gat);
  NR3 NOR3_60(n935gat,n938gat,n941gat,n942gat);
  NR3 NOR3_61(n936gat,n943gat,n939gat,n942gat);
  NR3 NOR3_62(n937gat,n943gat,n941gat,n940gat);
  NR2 NOR2_47(n746gat,n2716gat,n2723gat);
  NR2 NOR2_48(n360gat,n2859gat,n2727gat);
  NR3 NOR3_63(n710gat,n714gat,n715gat,n716gat);
  NR3 NOR3_64(n711gat,n714gat,n717gat,n718gat);
  NR3 NOR3_65(n712gat,n719gat,n715gat,n718gat);
  NR3 NOR3_66(n713gat,n719gat,n717gat,n716gat);
  NR3 NOR3_67(n729gat,n733gat,n734gat,n735gat);
  NR3 NOR3_68(n730gat,n733gat,n736gat,n737gat);
  NR3 NOR3_69(n731gat,n738gat,n734gat,n737gat);
  NR3 NOR3_70(n732gat,n738gat,n736gat,n735gat);
  NR3 NOR3_71(n494gat,n498gat,n499gat,n500gat);
  NR3 NOR3_72(n495gat,n498gat,n501gat,n502gat);
  NR3 NOR3_73(n496gat,n503gat,n499gat,n502gat);
  NR3 NOR3_74(n497gat,n503gat,n501gat,n500gat);
  NR3 NOR3_75(n505gat,n509gat,n510gat,n511gat);
  NR3 NOR3_76(n506gat,n509gat,n512gat,n513gat);
  NR3 NOR3_77(n507gat,n514gat,n510gat,n513gat);
  NR3 NOR3_78(n508gat,n514gat,n512gat,n511gat);
  NR4 NOR4_1(n564gat,n3029gat,n2863gat,n2855gat,n374gat);
  NR3 NOR3_79(n86gat,n743gat,n294gat,n17gat);
  NR2 NOR2_49(n78gat,n2784gat,n79gat);
  NR2 NOR2_50(n767gat,n219gat,n2731gat);
  NR2 NOR2_51(n286gat,n289gat,n2723gat);
  NR2 NOR2_52(n287gat,n289gat,n2715gat);
  NR2 NOR2_53(n288gat,n289gat,n2726gat);
  NR3 NOR3_80(n181gat,n286gat,n179gat,n188gat);
  NR2 NOR2_54(n182gat,n72gat,n2720gat);
  NR2 NOR2_55(n653gat,n2718gat,n111gat);
  NR2 NOR2_56(n867gat,n219gat,n2775gat);
  NR2 NOR2_57(n771gat,n2838gat,n111gat);
  NR2 NOR2_58(n964gat,n111gat,n2711gat);
  NR2 NOR2_59(n961gat,n219gat,n2734gat);
  NR3 NOR3_81(n804gat,n808gat,n809gat,n810gat);
  NR3 NOR3_82(n805gat,n808gat,n811gat,n812gat);
  NR3 NOR3_83(n806gat,n813gat,n809gat,n812gat);
  NR3 NOR3_84(n807gat,n813gat,n811gat,n810gat);
  NR3 NOR3_85(n587gat,n591gat,n592gat,n593gat);
  NR3 NOR3_86(n588gat,n591gat,n594gat,n595gat);
  NR3 NOR3_87(n589gat,n596gat,n592gat,n595gat);
  NR3 NOR3_88(n590gat,n596gat,n594gat,n593gat);
  NR2 NOR2_60(n447gat,n2836gat,n111gat);
  NR2 NOR2_61(n445gat,n2778gat,n219gat);
  NR3 NOR3_89(n687gat,n691gat,n692gat,n693gat);
  NR3 NOR3_90(n688gat,n691gat,n694gat,n695gat);
  NR3 NOR3_91(n689gat,n696gat,n692gat,n695gat);
  NR3 NOR3_92(n690gat,n696gat,n694gat,n693gat);
  NR3 NOR3_93(n568gat,n572gat,n573gat,n574gat);
  NR3 NOR3_94(n569gat,n572gat,n575gat,n576gat);
  NR3 NOR3_95(n570gat,n577gat,n573gat,n576gat);
  NR3 NOR3_96(n571gat,n577gat,n575gat,n574gat);
  NR3 NOR3_97(n187gat,n189gat,n287gat,n188gat);
  NR2 NOR2_62(n197gat,n194gat,n297gat);
  NR3 NOR3_98(n15gat,n637gat,n17gat,n293gat);
  NR2 NOR2_63(n22gat,n92gat,n21gat);
  NR2 NOR2_64(n93gat,n197gat,n22gat);
  NR2 NOR2_65(n769gat,n93gat,n2731gat);
  NR3 NOR3_99(n2534gat,n2624gat,n2489gat,n2621gat);
  NR3 NOR3_100(n2430gat,n2533gat,n2486gat,n2429gat);
  NR2 NOR2_66(n1606gat,n3020gat,n270gat);
  NR2 NOR2_67(n2239gat,n2850gat,n3019gat);
  NR3 NOR3_101(n1934gat,n2470gat,n1935gat,n2239gat);
  NR2 NOR2_68(n1610gat,n1698gat,n1543gat);
  NR2 NOR2_69(n1692gat,n1879gat,n1762gat);
  NR2 NOR2_70(n2433gat,n2432gat,n2154gat);
  NR3 NOR3_102(n2531gat,n2488gat,n2625gat,n2621gat);
  NR3 NOR3_103(n2480gat,n2530gat,n2482gat,n2486gat);
  NR2 NOR2_71(n2427gat,n2426gat,n2153gat);
  NR2 NOR2_72(n2428gat,n2433gat,n2427gat);
  NR2 NOR2_73(n1778gat,n3026gat,n1779gat);
  NR2 NOR2_74(n1609gat,n1503gat,n3025gat);
  NR2 NOR2_75(n1702gat,n3024gat,n1615gat);
  NR2 NOR2_76(n1700gat,n1701gat,n3023gat);
  NR4 NOR4_2(n1604gat,n1778gat,n1609gat,n1702gat,n1700gat);
  NR2 NOR2_77(n1076gat,n93gat,n2775gat);
  NR2 NOR2_78(n766gat,n93gat,n2734gat);
  NR3 NOR3_104(n1185gat,n1189gat,n1190gat,n1191gat);
  NR3 NOR3_105(n1186gat,n1189gat,n1192gat,n1193gat);
  NR3 NOR3_106(n1187gat,n1194gat,n1190gat,n1193gat);
  NR3 NOR3_107(n1188gat,n1194gat,n1192gat,n1191gat);
  NR2 NOR2_79(n645gat,n2792gat,n93gat);
  NR2 NOR2_80(n646gat,n93gat,n2669gat);
  NR2 NOR2_81(n1383gat,n1280gat,n1225gat);
  NR2 NOR2_82(n1327gat,n1281gat,n1224gat);
  NR2 NOR2_83(n651gat,n93gat,n2778gat);
  NR2 NOR2_84(n652gat,n2789gat,n93gat);
  NR2 NOR2_85(n765gat,n2781gat,n93gat);
  NR3 NOR3_108(n1202gat,n1206gat,n1207gat,n1208gat);
  NR3 NOR3_109(n1203gat,n1206gat,n1209gat,n1210gat);
  NR3 NOR3_110(n1204gat,n1211gat,n1207gat,n1210gat);
  NR3 NOR3_111(n1205gat,n1211gat,n1209gat,n1208gat);
  NR3 NOR3_112(n1270gat,n1274gat,n1275gat,n1276gat);
  NR3 NOR3_113(n1271gat,n1274gat,n1277gat,n1278gat);
  NR3 NOR3_114(n1272gat,n1279gat,n1275gat,n1278gat);
  NR3 NOR3_115(n1273gat,n1279gat,n1277gat,n1276gat);
  NR2 NOR2_86(n763gat,n2672gat,n93gat);
  NR2 NOR2_87(n1287gat,n1284gat,n1195gat);
  NR2 NOR2_88(n1285gat,n1196gat,n1269gat);
  NR2 NOR2_89(n853gat,n740gat,n2148gat);
  NR2 NOR2_90(n793gat,n2852gat,n851gat);
  NR2 NOR2_91(n854gat,n2148gat,n374gat);
  NR2 NOR2_92(n556gat,n2672gat,n852gat);
  NR2 NOR2_93(n795gat,n2731gat,n852gat);
  NR2 NOR2_94(n656gat,n851gat,n2718gat);
  NR2 NOR2_95(n794gat,n852gat,n2775gat);
  NR2 NOR2_96(n773gat,n851gat,n2838gat);
  NR2 NOR2_97(n965gat,n2711gat,n851gat);
  NR2 NOR2_98(n960gat,n2734gat,n852gat);
  NR3 NOR3_116(n780gat,n784gat,n785gat,n786gat);
  NR3 NOR3_117(n781gat,n784gat,n787gat,n788gat);
  NR3 NOR3_118(n782gat,n789gat,n785gat,n788gat);
  NR3 NOR3_119(n783gat,n789gat,n787gat,n786gat);
  NR2 NOR2_99(n555gat,n852gat,n2792gat);
  NR2 NOR2_100(n450gat,n851gat,n2846gat);
  NR2 NOR2_101(n654gat,n851gat,n2844gat);
  NR2 NOR2_102(n557gat,n2669gat,n852gat);
  NR2 NOR2_103(n874gat,n559gat,n365gat);
  NR2 NOR2_104(n132gat,n560gat,n364gat);
  NR2 NOR2_105(n649gat,n2778gat,n852gat);
  NR2 NOR2_106(n449gat,n2836gat,n851gat);
  NR2 NOR2_107(n791gat,n851gat,n2840gat);
  NR2 NOR2_108(n650gat,n852gat,n2789gat);
  NR2 NOR2_109(n774gat,n2842gat,n851gat);
  NR2 NOR2_110(n764gat,n852gat,n2781gat);
  NR3 NOR3_120(n222gat,n226gat,n227gat,n228gat);
  NR3 NOR3_121(n223gat,n226gat,n229gat,n230gat);
  NR3 NOR3_122(n224gat,n231gat,n227gat,n230gat);
  NR3 NOR3_123(n225gat,n231gat,n229gat,n228gat);
  NR3 NOR3_124(n121gat,n125gat,n126gat,n127gat);
  NR3 NOR3_125(n122gat,n125gat,n128gat,n129gat);
  NR3 NOR3_126(n123gat,n130gat,n126gat,n129gat);
  NR3 NOR3_127(n124gat,n130gat,n128gat,n127gat);
  NR2 NOR2_111(n2460gat,n666gat,n120gat);
  NR2 NOR2_112(n2423gat,n665gat,n1601gat);
  NR3 NOR3_128(n2594gat,n3017gat,n2520gat,n2597gat);
  NR3 NOR3_129(n2569gat,n2573gat,n2574gat,n2575gat);
  NR3 NOR3_130(n2570gat,n2573gat,n2576gat,n2577gat);
  NR3 NOR3_131(n2571gat,n2578gat,n2574gat,n2577gat);
  NR3 NOR3_132(n2572gat,n2578gat,n2576gat,n2575gat);
  NR3 NOR3_133(n2410gat,n2414gat,n2415gat,n2416gat);
  NR3 NOR3_134(n2411gat,n2414gat,n2417gat,n2418gat);
  NR3 NOR3_135(n2412gat,n2419gat,n2415gat,n2418gat);
  NR3 NOR3_136(n2413gat,n2419gat,n2417gat,n2416gat);
  NR2 NOR2_113(n2583gat,n2582gat,n2585gat);
  NR2 NOR2_114(n2580gat,n2582gat,n2583gat);
  NR2 NOR2_115(n2581gat,n2583gat,n2585gat);
  NR2 NOR2_116(n2567gat,n2493gat,n2388gat);
  NR2 NOR2_117(n2499gat,n2389gat,n2494gat);
  NR2 NOR2_118(n299gat,n2268gat,n2338gat);
  NR2 NOR2_119(n207gat,n2337gat,n2269gat);
  NR2 NOR2_120(n2650gat,n2649gat,n2652gat);
  NR2 NOR2_121(n2647gat,n2649gat,n2650gat);
  NR2 NOR2_122(n2648gat,n2650gat,n2652gat);
  NR3 NOR3_137(n2602gat,n2606gat,n2607gat,n2608gat);
  NR3 NOR3_138(n2603gat,n2606gat,n2609gat,n2610gat);
  NR3 NOR3_139(n2604gat,n2611gat,n2607gat,n2610gat);
  NR3 NOR3_140(n2605gat,n2611gat,n2609gat,n2608gat);
  NR3 NOR3_141(n2546gat,n2550gat,n2551gat,n2552gat);
  NR3 NOR3_142(n2547gat,n2550gat,n2553gat,n2554gat);
  NR3 NOR3_143(n2548gat,n2555gat,n2551gat,n2554gat);
  NR3 NOR3_144(n2549gat,n2555gat,n2553gat,n2552gat);
  NR2 NOR2_123(n2617gat,n2616gat,n2619gat);
  NR2 NOR2_124(n2614gat,n2616gat,n2617gat);
  NR2 NOR2_125(n2615gat,n2617gat,n2619gat);
  NR4 NOR4_3(n2655gat,n2508gat,n2656gat,n2500gat,n2504gat);
  NR3 NOR3_145(n2293gat,n2353gat,n2284gat,n2443gat);
  NR2 NOR2_126(n2219gat,n2354gat,n2214gat);
  NR2 NOR2_127(n1529gat,n1528gat,n1523gat);
  NR2 NOR2_128(n1704gat,n3027gat,n1706gat);
  NR2 NOR2_129(n2461gat,n120gat,n2666gat);
  NR2 NOR2_130(n2421gat,n1601gat,n1704gat);
  NR2 NOR2_131(n1598gat,n1592gat,n2422gat);
  NR2 NOR2_132(n2218gat,n2214gat,n2290gat);
  NR3 NOR3_146(n2358gat,n2285gat,n2356gat,n2355gat);
  NR2 NOR2_133(n1415gat,n2081gat,n2359gat);
  NR2 NOR2_134(n1153gat,n1414gat,n566gat);
  NR3 NOR3_147(n2292gat,n2443gat,n2284gat,n2285gat);
  NR2 NOR2_135(n1416gat,n2081gat,n1480gat);
  NR2 NOR2_136(n1151gat,n1301gat,n1150gat);
  NR3 NOR3_148(n2306gat,n2356gat,n2284gat,n2285gat);
  NR2 NOR2_137(n1481gat,n2081gat,n2011gat);
  NR2 NOR2_138(n982gat,n873gat,n1478gat);
  NR3 NOR3_149(n2357gat,n2285gat,n2355gat,n2443gat);
  NR2 NOR2_139(n1347gat,n2081gat,n1410gat);
  NR2 NOR2_140(n877gat,n875gat,n876gat);
  NR2 NOR2_141(n1484gat,n2081gat,n1528gat);
  NR2 NOR2_142(n1159gat,n1160gat,n1084gat);
  NR3 NOR3_150(n2363gat,n2353gat,n2356gat,n2355gat);
  NR2 NOR2_143(n1483gat,n2081gat,n1482gat);
  NR2 NOR2_144(n1158gat,n983gat,n1157gat);
  NR3 NOR3_151(n2364gat,n2353gat,n2284gat,n2356gat);
  NR2 NOR2_145(n1308gat,n2081gat,n1530gat);
  NR2 NOR2_146(n1156gat,n985gat,n1307gat);
  NR3 NOR3_152(n2291gat,n2353gat,n2355gat,n2443gat);
  NR2 NOR2_147(n1349gat,n1479gat,n2081gat);
  NR2 NOR2_148(n1155gat,n1085gat,n1348gat);
  NR3 NOR3_153(n1154gat,n1598gat,n2930gat,n2957gat);
  NR2 NOR2_149(n1703gat,n1705gat,n3028gat);
  NR2 NOR2_150(n1608gat,n1704gat,n1703gat);
  NR2 NOR2_151(n1411gat,n1154gat,n1608gat);
  NR2 NOR2_152(n2223gat,n2354gat,n2217gat);
  NR2 NOR2_153(n1438gat,n1591gat,n1480gat);
  NR2 NOR2_154(n1625gat,n3021gat,n1628gat);
  NR2 NOR2_155(n1626gat,n1627gat,n3022gat);
  NR3 NOR3_154(n1831gat,n1832gat,n1765gat,n1878gat);
  NR2 NOR2_156(n1443gat,n1442gat,n706gat);
  NR2 NOR2_157(n1325gat,n1444gat,n164gat);
  NR2 NOR2_158(n1441gat,n1437gat,n1378gat);
  NR2 NOR2_159(n1321gat,n1442gat,n837gat);
  NR2 NOR2_160(n1320gat,n1444gat,n278gat);
  NR2 NOR2_161(n1486gat,n1482gat,n1591gat);
  NR2 NOR2_162(n1440gat,n1322gat,n1439gat);
  NR2 NOR2_163(n1426gat,n2011gat,n1591gat);
  NR2 NOR2_164(n1368gat,n1442gat,n613gat);
  NR2 NOR2_165(n1258gat,n274gat,n1444gat);
  NR2 NOR2_166(n1371gat,n1370gat,n1369gat);
  NR2 NOR2_167(n1365gat,n1479gat,n1591gat);
  NR2 NOR2_168(n1373gat,n833gat,n1442gat);
  NR2 NOR2_169(n1372gat,n282gat,n1444gat);
  NR2 NOR2_170(n1367gat,n1366gat,n1374gat);
  NR2 NOR2_171(n2220gat,n2290gat,n2217gat);
  NR2 NOR2_172(n1423gat,n2162gat,n1530gat);
  NR2 NOR2_173(n1498gat,n1609gat,n1427gat);
  NR2 NOR2_174(n1504gat,n1450gat,n1498gat);
  NR2 NOR2_175(n1607gat,n2082gat,n1609gat);
  NR2 NOR2_176(n1494gat,n1528gat,n2162gat);
  NR2 NOR2_177(n1502gat,n1607gat,n1449gat);
  NR2 NOR2_178(n1250gat,n1603gat,n815gat);
  NR2 NOR2_179(n1103gat,n956gat,n1590gat);
  NR2 NOR2_180(n1417gat,n2162gat,n1480gat);
  NR2 NOR2_181(n1352gat,n1248gat,n1418gat);
  NR2 NOR2_182(n1304gat,n1590gat,n1067gat);
  NR2 NOR2_183(n1249gat,n679gat,n1603gat);
  NR2 NOR2_184(n1419gat,n2162gat,n1479gat);
  NR2 NOR2_185(n1351gat,n1306gat,n1353gat);
  NR2 NOR2_186(n1246gat,n864gat,n1590gat);
  NR2 NOR2_187(n1161gat,n583gat,n1603gat);
  NR2 NOR2_188(n1422gat,n2011gat,n2162gat);
  NR2 NOR2_189(n1303gat,n1247gat,n1355gat);
  NR2 NOR2_190(n1291gat,n1603gat,n579gat);
  NR2 NOR2_191(n1245gat,n1590gat,n860gat);
  NR2 NOR2_192(n1485gat,n1482gat,n2162gat);
  NR2 NOR2_193(n1302gat,n1300gat,n1487gat);
  NR2 NOR2_194(n1163gat,n882gat,n1603gat);
  NR2 NOR2_195(n1102gat,n1297gat,n1590gat);
  NR2 NOR2_196(n1354gat,n1591gat,n1530gat);
  NR2 NOR2_197(n1360gat,n1164gat,n1356gat);
  NR2 NOR2_198(n1435gat,n1591gat,n1528gat);
  NR2 NOR2_199(n1101gat,n1590gat,n1293gat);
  NR2 NOR2_200(n996gat,n1603gat,n823gat);
  NR2 NOR2_201(n1359gat,n1436gat,n1106gat);
  NR2 NOR2_202(n1421gat,n2162gat,n2359gat);
  NR2 NOR2_203(n1104gat,n1079gat,n1590gat);
  NR2 NOR2_204(n887gat,n1603gat,n683gat);
  NR2 NOR2_205(n1358gat,n1425gat,n1105gat);
  NR2 NOR2_206(n1420gat,n1410gat,n2162gat);
  NR2 NOR2_207(n1305gat,n1147gat,n1590gat);
  NR2 NOR2_208(n1162gat,n698gat,n1603gat);
  NR2 NOR2_209(n1357gat,n1424gat,n1309gat);
  NR4 NOR4_4(n1428gat,n2978gat,n2982gat,n2973gat,n2977gat);
  NR2 NOR2_210(n1794gat,n1673gat,n1719gat);
  NR2 NOR2_211(n1796gat,n1858gat,n1635gat);
  NR2 NOR2_212(n1792gat,n1794gat,n1796gat);
  NR3 NOR3_155(n1865gat,n1989gat,n1918gat,n1986gat);
  NR3 NOR3_156(n1861gat,n1866gat,n2216gat,n1988gat);
  NR2 NOR2_213(n1793gat,n1792gat,n1735gat);
  NR2 NOR2_214(n1406gat,n1428gat,n1387gat);
  NR3 NOR3_157(n1780gat,n1777gat,n1625gat,n1626gat);
  NR2 NOR2_215(n2016gat,n2019gat,n1878gat);
  NR2 NOR2_216(n2664gat,n2850gat,n3018gat);
  NR3 NOR3_158(n1666gat,n1986gat,n2212gat,n1991gat);
  NR3 NOR3_159(n1578gat,n2152gat,n2351gat,n1665gat);
  NR2 NOR2_217(n1516gat,n1551gat,n1517gat);
  NR3 NOR3_160(n1864gat,n1858gat,n1495gat,n2090gat);
  NR2 NOR2_218(n1565gat,n1735gat,n1552gat);
  NR2 NOR2_219(n1921gat,n1738gat,n1673gat);
  NR2 NOR2_220(n1798gat,n1739gat,n1673gat);
  NR3 NOR3_161(n1920gat,n1864gat,n1921gat,n1798gat);
  NR2 NOR2_221(n1926gat,n1925gat,n1635gat);
  NR2 NOR2_222(n1916gat,n1917gat,n1859gat);
  NR2 NOR2_223(n1994gat,n1719gat,n1922gat);
  NR2 NOR2_224(n1924gat,n1743gat,n1923gat);
  NR4 NOR4_5(n2078gat,n1926gat,n1916gat,n1994gat,n1924gat);
  NR2 NOR2_225(n1690gat,n1700gat,n1702gat);
  NR3 NOR3_162(n1660gat,n1918gat,n1986gat,n2212gat);
  NR3 NOR3_163(n1576gat,n2351gat,n1988gat,n1661gat);
  NR2 NOR2_226(n1733gat,n1673gat,n1572gat);
  NR3 NOR3_164(n1582gat,n2283gat,n1991gat,n2212gat);
  NR3 NOR3_165(n1577gat,n1520gat,n2351gat,n1988gat);
  NR2 NOR2_227(n1581gat,n1858gat,n1580gat);
  NR3 NOR3_166(n2129gat,n2189gat,n2134gat,n2261gat);
  NR4 NOR4_6(n2079gat,n2078gat,n2178gat,n1990gat,n2128gat);
  NR4 NOR4_7(n1695gat,n1609gat,n1778gat,n1704gat,n1703gat);
  NR3 NOR3_167(n2073gat,n2078gat,n1990gat,n2181gat);
  NR2 NOR2_228(n1696gat,n1707gat,n1698gat);
  NR2 NOR2_229(n1758gat,n1311gat,n1773gat);
  NR3 NOR3_168(n1574gat,n1719gat,n1673gat,n1444gat);
  NR3 NOR3_169(n1573gat,n1444gat,n1858gat,n1635gat);
  NR2 NOR2_230(n1521gat,n2283gat,n1991gat);
  NR2 NOR2_231(n1737gat,n2212gat,n2152gat);
  NR3 NOR3_170(n1732gat,n1515gat,n1736gat,n1658gat);
  NR3 NOR3_171(n1723gat,n1659gat,n1722gat,n1724gat);
  NR2 NOR2_232(n1663gat,n1986gat,n1918gat);
  NR3 NOR3_172(n1655gat,n1736gat,n1662gat,n1658gat);
  NR3 NOR3_173(n1647gat,n1656gat,n1659gat,n1554gat);
  NR2 NOR2_233(n1667gat,n1991gat,n1986gat);
  NR3 NOR3_174(n1570gat,n1736gat,n1658gat,n1670gat);
  NR3 NOR3_175(n1646gat,n1569gat,n1659gat,n1566gat);
  NR2 NOR2_234(n1575gat,n1918gat,n2283gat);
  NR3 NOR3_176(n1728gat,n1568gat,n1736gat,n1658gat);
  NR3 NOR3_177(n1650gat,n1727gat,n1659gat,n1640gat);
  NR2 NOR2_235(n1801gat,n2152gat,n1989gat);
  NR3 NOR3_178(n1731gat,n1658gat,n1515gat,n1797gat);
  NR3 NOR3_179(n1649gat,n1560gat,n1659gat,n1730gat);
  NR3 NOR3_180(n1571gat,n1670gat,n1658gat,n1797gat);
  NR3 NOR3_181(n1563gat,n1561gat,n1562gat,n1659gat);
  NR2 NOR2_236(n1734gat,n1988gat,n2212gat);
  NR3 NOR3_182(n1669gat,n1668gat,n1742gat,n1670gat);
  NR2 NOR2_237(n1654gat,n1671gat,n1659gat);
  NR3 NOR3_183(n1657gat,n1662gat,n1797gat,n1658gat);
  NR3 NOR3_184(n1653gat,n1651gat,n1652gat,n1659gat);
  NR3 NOR3_185(n1729gat,n1658gat,n1797gat,n1568gat);
  NR3 NOR3_186(n1644gat,n1643gat,n1648gat,n1659gat);
  NR3 NOR3_187(n1726gat,n2992gat,n2986gat,n2991gat);
  NR2 NOR2_238(n1929gat,n1758gat,n1790gat);
  NR3 NOR3_188(n2009gat,n2016gat,n2664gat,n2004gat);
  NR3 NOR3_189(n1413gat,n1869gat,n672gat,n2591gat);
  NR2 NOR2_239(n1636gat,n1584gat,n1718gat);
  NR2 NOR2_240(n1401gat,n1584gat,n1590gat);
  NR3 NOR3_190(n1408gat,n1507gat,n1396gat,n1393gat);
  NR2 NOR2_241(n1476gat,n1858gat,n1590gat);
  NR3 NOR3_191(n1407gat,n1393gat,n1409gat,n1677gat);
  NR3 NOR3_192(n1412gat,n1411gat,n1406gat,n2981gat);
  NR3 NOR3_193(n2663gat,n2586gat,n2660gat,n2307gat);
  NR2 NOR2_242(n2662gat,n2660gat,n2586gat);
  NR2 NOR2_243(n2238gat,n2448gat,n2444gat);
  NR3 NOR3_194(n87gat,n743gat,n17gat,n293gat);
  NR2 NOR2_244(n200gat,n199gat,n92gat);
  NR3 NOR3_195(n184gat,n189gat,n188gat,n179gat);
  NR2 NOR2_245(n196gat,n297gat,n195gat);
  NR2 NOR2_246(n204gat,n200gat,n196gat);
  NR4 NOR4_8(n2163gat,n1790gat,n1310gat,n2664gat,n2168gat);
  NR2 NOR2_247(n2258gat,n2260gat,n2189gat);
  NR2 NOR2_248(n2255gat,n2261gat,n2188gat);
  NR3 NOR3_196(n2015gat,n2039gat,n1774gat,n1315gat);
  NR2 NOR2_249(n2017gat,n1790gat,n2016gat);
  NR2 NOR2_250(n2018gat,n2016gat,n2097gat);
  NR4 NOR4_9(n2014gat,n2035gat,n2093gat,n2018gat,n2664gat);
  NR2 NOR2_251(n2194gat,n2187gat,n1855gat);
  NR2 NOR2_252(n2192gat,n2184gat,n1855gat);
  NR2 NOR2_253(n2185gat,n2261gat,n2189gat);
  NR2 NOR2_254(n2132gat,n2133gat,n2131gat);
  NR2 NOR2_255(n2130gat,n2134gat,n2185gat);
  NR2 NOR2_256(n2057gat,n2049gat,n1855gat);
  NR2 NOR2_257(n2250gat,n2248gat,n2264gat);
  NR2 NOR2_258(n2249gat,n2265gat,n3006gat);
  NR2 NOR2_259(n2329gat,n1855gat,n3007gat);
  NR2 NOR2_260(n1958gat,n1963gat,n1886gat);
  NR3 NOR3_197(n1895gat,n1845gat,n1891gat,n1968gat);
  NR2 NOR2_261(n1710gat,n1709gat,n1629gat);
  NR2 NOR2_262(n1630gat,n1895gat,n1631gat);
  NR2 NOR2_263(n2195gat,n2200gat,n1855gat);
  NR2 NOR2_264(n2556gat,n1711gat,n2437gat);
  NR2 NOR2_265(n2539gat,n2048gat,n2437gat);
  NR3 NOR3_198(n1894gat,n1968gat,n1891gat,n1969gat);
  NR2 NOR2_266(n1847gat,n1958gat,n1845gat);
  NR2 NOR2_267(n1846gat,n1845gat,n1893gat);
  NR2 NOR2_268(n2436gat,n2437gat,n1892gat);
  NR2 NOR2_269(n2055gat,n1891gat,n1958gat);
  NR2 NOR2_270(n1967gat,n1893gat,n1968gat);
  NR2 NOR2_271(n2387gat,n2056gat,n2437gat);
  NR2 NOR2_272(n1959gat,n1956gat,n1963gat);
  NR2 NOR2_273(n1957gat,n1886gat,n1887gat);
  NR2 NOR2_274(n2330gat,n2437gat,n1961gat);
  NR2 NOR2_275(n2147gat,n2988gat,n1855gat);
  NR2 NOR2_276(n2498gat,n2199gat,n2328gat);
  NR2 NOR2_277(n2193gat,n2393gat,n2439gat);
  NR2 NOR2_278(n2211gat,n2193gat,n2402gat);
  NR2 NOR2_279(n2210gat,n2401gat,n2151gat);
  NR2 NOR2_280(n2396gat,n2199gat,n2209gat);
  NR2 NOR2_281(n2053gat,n2393gat,n2438gat);
  NR2 NOR2_282(n1964gat,n2392gat,n2439gat);
  NR2 NOR2_283(n2198gat,n2199gat,n2058gat);
  NR3 NOR3_199(n2215gat,n2346gat,n2151gat,n2402gat);
  NR2 NOR2_284(n2350gat,n2405gat,n2349gat);
  NR2 NOR2_285(n2282gat,n2406gat,n2215gat);
  NR2 NOR2_286(n2197gat,n2199gat,n2281gat);
  NR3 NOR3_200(n2213gat,n2402gat,n2151gat,n2345gat);
  NR2 NOR2_287(n2150gat,n2401gat,n2346gat);
  NR2 NOR2_288(n2149gat,n2193gat,n2346gat);
  NR2 NOR2_289(n2196gat,n2199gat,n2146gat);
  NR3 NOR3_201(n1882gat,n2124gat,n2115gat,n2239gat);
  NR2 NOR2_290(n1962gat,n1963gat,n1893gat);
  NR2 NOR2_291(n1896gat,n2995gat,n1895gat);
  NR2 NOR2_292(n1972gat,n1974gat,n1970gat);
  NR2 NOR2_293(n1971gat,n1896gat,n1973gat);
  NR2 NOR2_294(n2559gat,n2999gat,n2437gat);
  NR2 NOR2_295(n2331gat,n2393gat,n2401gat);
  NR2 NOR2_296(n2352gat,n3011gat,n2215gat);
  NR2 NOR2_297(n2566gat,n2643gat,n2564gat);
  NR2 NOR2_298(n2565gat,n2352gat,n2642gat);
  NR2 NOR2_299(n2637gat,n3015gat,n2199gat);
  NR3 NOR3_202(n84gat,n296gat,n17gat,n294gat);
  NR2 NOR2_300(n89gat,n88gat,n2784gat);
  NR2 NOR2_301(n110gat,n182gat,n89gat);
  NR2 NOR2_302(n1074gat,n2775gat,n110gat);
  NR3 NOR3_203(n141gat,n155gat,n253gat,n150gat);
  NR2 NOR2_303(n38gat,n151gat,n233gat);
  NR2 NOR2_304(n37gat,n151gat,n154gat);
  NR2 NOR2_305(n872gat,n375gat,n800gat);
  NR2 NOR2_306(n234gat,n155gat,n233gat);
  NR2 NOR2_307(n137gat,n154gat,n253gat);
  NR2 NOR2_308(n378gat,n375gat,n235gat);
  NR2 NOR2_309(n377gat,n110gat,n2778gat);
  NR2 NOR2_310(n869gat,n219gat,n2792gat);
  NR2 NOR2_311(n212gat,n182gat,n78gat);
  NR3 NOR3_204(n250gat,n329gat,n387gat,n334gat);
  NR2 NOR2_312(n249gat,n386gat,n330gat);
  NR2 NOR2_313(n248gat,n330gat,n1490gat);
  NR2 NOR2_314(n453gat,n372gat,n452gat);
  NR2 NOR2_315(n448gat,n111gat,n2846gat);
  NR2 NOR2_316(n974gat,n2844gat,n111gat);
  NR2 NOR2_317(n251gat,n1490gat,n387gat);
  NR2 NOR2_318(n244gat,n334gat,n386gat);
  NR2 NOR2_319(n973gat,n372gat,n333gat);
  NR2 NOR2_320(n870gat,n2669gat,n219gat);
  NR2 NOR2_321(n975gat,n111gat,n2852gat);
  NR3 NOR3_205(n246gat,n330gat,n325gat,n334gat);
  NR2 NOR2_322(n245gat,n386gat,n334gat);
  NR2 NOR2_323(n460gat,n462gat,n2884gat);
  NR2 NOR2_324(n459gat,n457gat,n461gat);
  NR2 NOR2_325(n972gat,n372gat,n458gat);
  NR2 NOR2_326(n969gat,n219gat,n2672gat);
  NR2 NOR2_327(n971gat,n111gat,n2840gat);
  NR3 NOR3_206(n247gat,n334gat,n387gat,n330gat);
  NR2 NOR2_328(n145gat,n144gat,n325gat);
  NR2 NOR2_329(n143gat,n326gat,n247gat);
  NR2 NOR2_330(n970gat,n372gat,n878gat);
  NR2 NOR2_331(n968gat,n2789gat,n219gat);
  NR2 NOR2_332(n772gat,n111gat,n2842gat);
  NR3 NOR3_207(n142gat,n382gat,n326gat,n144gat);
  NR2 NOR2_333(n40gat,n325gat,n383gat);
  NR2 NOR2_334(n39gat,n383gat,n247gat);
  NR2 NOR2_335(n451gat,n134gat,n372gat);
  NR2 NOR2_336(n446gat,n219gat,n2781gat);
  NR3 NOR3_208(n139gat,n253gat,n151gat,n254gat);
  NR2 NOR2_337(n136gat,n253gat,n154gat);
  NR2 NOR2_338(n391gat,n252gat,n468gat);
  NR2 NOR2_339(n390gat,n469gat,n2877gat);
  NR2 NOR2_340(n1083gat,n381gat,n375gat);
  NR2 NOR2_341(n1077gat,n110gat,n2672gat);
  NR3 NOR3_209(n140gat,n151gat,n253gat,n155gat);
  NR2 NOR2_342(n242gat,n254gat,n241gat);
  NR2 NOR2_343(n240gat,n255gat,n140gat);
  NR2 NOR2_344(n871gat,n802gat,n375gat);
  NR2 NOR2_345(n797gat,n110gat,n2734gat);
  NR3 NOR3_210(n324gat,n255gat,n146gat,n241gat);
  NR2 NOR2_346(n238gat,n147gat,n254gat);
  NR2 NOR2_347(n237gat,n140gat,n147gat);
  NR2 NOR2_348(n1082gat,n375gat,n380gat);
  NR2 NOR2_349(n796gat,n2731gat,n110gat);
  NR3 NOR3_211(n85gat,n17gat,n294gat,n637gat);
  NR3 NOR3_212(n180gat,n286gat,n188gat,n287gat);
  NR2 NOR2_350(n68gat,n85gat,n180gat);
  NR3 NOR3_213(n186gat,n189gat,n287gat,n288gat);
  NR2 NOR2_351(n357gat,n2726gat,n2860gat);
  NR3 NOR3_214(n82gat,n16gat,n295gat,n637gat);
  NR2 NOR2_352(n12gat,n186gat,n82gat);
  NR2 NOR2_353(n1599gat,n1691gat,n336gat);
  NR2 NOR2_354(n1613gat,n1544gat,n1698gat);
  NR3 NOR3_215(n1756gat,n2512gat,n1769gat,n1773gat);
  NR2 NOR2_355(n1586gat,n1869gat,n1683gat);
  NR3 NOR3_216(n1755gat,n1769gat,n1773gat,n2512gat);
  NR3 NOR3_217(n2538gat,n2620gat,n2625gat,n2488gat);
  NR3 NOR3_218(n2483gat,n2537gat,n2482gat,n2486gat);
  NR2 NOR2_356(n1391gat,n1513gat,n2442gat);
  NR3 NOR3_219(n1471gat,n1334gat,n1858gat,n1604gat);
  NR2 NOR2_357(n1469gat,n1858gat,n1608gat);
  NR3 NOR3_220(n1472gat,n1476gat,n1471gat,n1469gat);
  NR2 NOR2_358(n1927gat,n1790gat,n1635gat);
  NR2 NOR2_359(n1470gat,n1472gat,n1747gat);
  NR3 NOR3_221(n1402gat,n1858gat,n1393gat,n1604gat);
  NR2 NOR2_360(n1400gat,n1674gat,n1403gat);
  NR2 NOR2_361(n1567gat,n1634gat,n1735gat);
  NR3 NOR3_222(n1399gat,n1806gat,n1338gat,n1584gat);
  NR4 NOR4_10(n1564gat,n1584gat,n1719gat,n1790gat,n1576gat);
  NR2 NOR2_362(n1600gat,n1685gat,n1427gat);
  NR3 NOR3_223(n1519gat,n1584gat,n1339gat,n1600gat);
  NR2 NOR2_363(n1397gat,n1519gat,n1401gat);
  NR2 NOR2_364(n1398gat,n1455gat,n1397gat);
  NR2 NOR2_365(n2008gat,n2012gat,n1774gat);
  NR2 NOR2_366(n2005gat,n2002gat,n2857gat);
  NR2 NOR2_367(n1818gat,n1823gat,n2005gat);
  NR3 NOR3_224(n1759gat,n1818gat,n1935gat,n2765gat);
  NR3 NOR3_225(n1686gat,n1774gat,n1869gat,n1684gat);
  NR2 NOR2_368(n1533gat,n1524gat,n1403gat);
  NR3 NOR3_226(n1863gat,n1991gat,n2283gat,n1989gat);
  NR3 NOR3_227(n1860gat,n1988gat,n2216gat,n1862gat);
  NR2 NOR2_369(n1915gat,n1859gat,n1919gat);
  NR2 NOR2_370(n1510gat,n1584gat,n1460gat);
  NR2 NOR2_371(n1800gat,n1635gat,n1919gat);
  NR2 NOR2_372(n1459gat,n1595gat,n1454gat);
  NR2 NOR2_373(n1458gat,n1510gat,n1459gat);
  NR2 NOR2_374(n1532gat,n1677gat,n1458gat);
  NR2 NOR2_375(n1467gat,n2289gat,n1468gat);
  NR3 NOR3_228(n1466gat,n1392gat,n1461gat,n1396gat);
  NR2 NOR2_376(n1531gat,n1507gat,n1477gat);
  NR2 NOR2_377(n1593gat,n1551gat,n1310gat);
  NR3 NOR3_229(n1602gat,n1594gat,n1587gat,n2989gat);
  NR3 NOR3_230(n1761gat,n2985gat,n1602gat,n1681gat);
  NR3 NOR3_231(n1760gat,n1681gat,n1602gat,n2985gat);
  NR3 NOR3_232(n1721gat,n2442gat,n1690gat,n1978gat);
  NR2 NOR2_378(n520gat,n374gat,n2862gat);
  NR2 NOR2_379(n519gat,n2854gat,n374gat);
  NR2 NOR2_380(n518gat,n520gat,n519gat);
  NR2 NOR2_381(n418gat,n374gat,n2723gat);
  NR2 NOR2_382(n411gat,n374gat,n2726gat);
  NR2 NOR2_383(n522gat,n374gat,n2859gat);
  NR2 NOR2_384(n516gat,n374gat,n2715gat);
  NR4 NOR4_11(n410gat,n417gat,n413gat,n412gat,n406gat);
  NR2 NOR2_385(n354gat,n411gat,n522gat);
  NR3 NOR3_233(n355gat,n517gat,n410gat,n354gat);
  NR2 NOR2_386(n408gat,n516gat,n407gat);
  NR2 NOR2_387(n526gat,n2859gat,n740gat);
  NR2 NOR2_388(n531gat,n740gat,n2854gat);
  NR2 NOR2_389(n530gat,n2862gat,n740gat);
  NR3 NOR3_234(n525gat,n526gat,n531gat,n530gat);
  NR2 NOR2_390(n356gat,n2726gat,n740gat);
  NR2 NOR2_391(n415gat,n2723gat,n740gat);
  NR2 NOR2_392(n521gat,n740gat,n2715gat);
  NR3 NOR3_235(n532gat,n527gat,n416gat,n528gat);
  NR2 NOR2_393(n359gat,n290gat,n358gat);
  NR2 NOR2_394(n420gat,n408gat,n359gat);
  NR2 NOR2_395(n523gat,n522gat,n356gat);
  NR2 NOR2_396(n634gat,n418gat,n521gat);
  NR2 NOR2_397(n414gat,n411gat,n415gat);
  NR3 NOR3_236(n635gat,n639gat,n634gat,n414gat);
  NR2 NOR2_398(n1100gat,n1297gat,n1111gat);
  NR3 NOR3_237(n630gat,n634gat,n523gat,n524gat);
  NR2 NOR2_399(n994gat,n1112gat,n882gat);
  NR3 NOR3_238(n629gat,n414gat,n634gat,n523gat);
  NR2 NOR2_400(n989gat,n721gat,n741gat);
  NR3 NOR3_239(n632gat,n414gat,n523gat,n633gat);
  NR2 NOR2_401(n880gat,n926gat,n566gat);
  NR3 NOR3_240(n636gat,n414gat,n633gat,n639gat);
  NR2 NOR2_402(n801gat,n672gat,n670gat);
  NR2 NOR2_403(n879gat,n2931gat,n801gat);
  NR2 NOR2_404(n1003gat,n420gat,n879gat);
  NR2 NOR2_405(n1255gat,n1123gat,n1225gat);
  NR2 NOR2_406(n1012gat,n1007gat,n918gat);
  NR2 NOR2_407(n905gat,n625gat,n1006gat);
  NR2 NOR2_408(n1009gat,n1255gat,n2943gat);
  NR2 NOR2_409(n409gat,n406gat,n407gat);
  NR2 NOR2_410(n292gat,n415gat,n356gat);
  NR2 NOR2_411(n291gat,n290gat,n292gat);
  NR2 NOR2_412(n419gat,n409gat,n291gat);
  NR2 NOR2_413(n902gat,n1009gat,n419gat);
  NR2 NOR2_414(n1099gat,n1111gat,n1293gat);
  NR2 NOR2_415(n998gat,n725gat,n741gat);
  NR2 NOR2_416(n995gat,n823gat,n1112gat);
  NR2 NOR2_417(n980gat,n875gat,n926gat);
  NR2 NOR2_418(n1001gat,n420gat,n1002gat);
  NR2 NOR2_419(n1175gat,n621gat,n1006gat);
  NR2 NOR2_420(n1174gat,n845gat,n1007gat);
  NR2 NOR2_421(n1243gat,n1281gat,n1123gat);
  NR2 NOR2_422(n1171gat,n2960gat,n1243gat);
  NR2 NOR2_423(n999gat,n419gat,n1171gat);
  NR2 NOR2_424(n1244gat,n1123gat,n1134gat);
  NR2 NOR2_425(n1323gat,n1007gat,n401gat);
  NR2 NOR2_426(n1264gat,n1006gat,n617gat);
  NR2 NOR2_427(n1265gat,n1244gat,n2969gat);
  NR2 NOR2_428(n892gat,n419gat,n1265gat);
  NR2 NOR2_429(n981gat,n926gat,n873gat);
  NR2 NOR2_430(n890gat,n741gat,n702gat);
  NR2 NOR2_431(n889gat,n1111gat,n1079gat);
  NR2 NOR2_432(n886gat,n683gat,n1112gat);
  NR2 NOR2_433(n891gat,n420gat,n888gat);
  NR2 NOR2_434(n904gat,n1006gat,n490gat);
  NR2 NOR2_435(n903gat,n1007gat,n397gat);
  NR2 NOR2_436(n1254gat,n1123gat,n1044gat);
  NR2 NOR2_437(n1008gat,n2942gat,n1254gat);
  NR2 NOR2_438(n900gat,n419gat,n1008gat);
  NR2 NOR2_439(n1152gat,n926gat,n1150gat);
  NR2 NOR2_440(n1092gat,n1147gat,n1111gat);
  NR2 NOR2_441(n997gat,n741gat,n393gat);
  NR2 NOR2_442(n993gat,n1112gat,n698gat);
  NR2 NOR2_443(n895gat,n420gat,n898gat);
  NR2 NOR2_444(n1094gat,n1112gat,n583gat);
  NR2 NOR2_445(n1093gat,n1111gat,n864gat);
  NR2 NOR2_446(n988gat,n340gat,n741gat);
  NR2 NOR2_447(n984gat,n926gat,n983gat);
  NR2 NOR2_448(n1178gat,n420gat,n1179gat);
  NR2 NOR2_449(n1267gat,n613gat,n1006gat);
  NR2 NOR2_450(n1257gat,n1007gat,n274gat);
  NR2 NOR2_451(n1253gat,n930gat,n1123gat);
  NR2 NOR2_452(n1266gat,n2965gat,n1253gat);
  NR2 NOR2_453(n1116gat,n419gat,n1266gat);
  NR2 NOR2_454(n1375gat,n1006gat,n706gat);
  NR2 NOR2_455(n1324gat,n164gat,n1007gat);
  NR2 NOR2_456(n1200gat,n1120gat,n1123gat);
  NR2 NOR2_457(n1172gat,n2961gat,n1200gat);
  NR2 NOR2_458(n899gat,n419gat,n1172gat);
  NR2 NOR2_459(n1091gat,n1111gat,n956gat);
  NR2 NOR2_460(n1088gat,n1085gat,n926gat);
  NR2 NOR2_461(n992gat,n815gat,n1112gat);
  NR2 NOR2_462(n987gat,n741gat,n159gat);
  NR2 NOR2_463(n896gat,n897gat,n420gat);
  NR2 NOR2_464(n1262gat,n837gat,n1006gat);
  NR2 NOR2_465(n1260gat,n1007gat,n278gat);
  NR2 NOR2_466(n1251gat,n1123gat,n1071gat);
  NR2 NOR2_467(n1259gat,n2967gat,n1251gat);
  NR2 NOR2_468(n901gat,n419gat,n1259gat);
  NR2 NOR2_469(n1098gat,n336gat,n741gat);
  NR2 NOR2_470(n1090gat,n1111gat,n860gat);
  NR2 NOR2_471(n986gat,n985gat,n926gat);
  NR2 NOR2_472(n885gat,n579gat,n1112gat);
  NR2 NOR2_473(n893gat,n894gat,n420gat);
  NR2 NOR2_474(n1097gat,n270gat,n741gat);
  NR2 NOR2_475(n1089gat,n1067gat,n1111gat);
  NR2 NOR2_476(n1087gat,n926gat,n1084gat);
  NR2 NOR2_477(n991gat,n1112gat,n679gat);
  NR2 NOR2_478(n1177gat,n1180gat,n420gat);
  NR2 NOR2_479(n1212gat,n1123gat,n1034gat);
  NR2 NOR2_480(n1326gat,n1007gat,n282gat);
  NR2 NOR2_481(n1261gat,n833gat,n1006gat);
  NR2 NOR2_482(n1263gat,n1212gat,n2968gat);
  NR2 NOR2_483(n1115gat,n1263gat,n419gat);
  NR2 NOR2_484(n977gat,n670gat,n671gat);
  NR3 NOR3_241(n631gat,n523gat,n633gat,n524gat);
  NR2 NOR2_485(n1096gat,n819gat,n1112gat);
  NR2 NOR2_486(n1095gat,n1240gat,n1111gat);
  NR2 NOR2_487(n990gat,n841gat,n741gat);
  NR2 NOR2_488(n979gat,n1601gat,n926gat);
  NR2 NOR2_489(n978gat,n2944gat,n2945gat);
  NR2 NOR2_490(n1004gat,n978gat,n420gat);
  NR2 NOR2_491(n1199gat,n1123gat,n1284gat);
  NR2 NOR2_492(n1176gat,n829gat,n1006gat);
  NR2 NOR2_493(n1173gat,n1007gat,n1025gat);
  NR2 NOR2_494(n1252gat,n1199gat,n2962gat);
  NR2 NOR2_495(n1000gat,n419gat,n1252gat);
  NR2 NOR2_496(n1029gat,n978gat,n455gat);
  NR2 NOR2_497(n1028gat,n455gat,n879gat);
  NR2 NOR2_498(n1031gat,n1002gat,n455gat);
  NR2 NOR2_499(n1030gat,n455gat,n888gat);
  NR2 NOR2_500(n1011gat,n455gat,n898gat);
  NR2 NOR2_501(n1181gat,n455gat,n1179gat);
  NR2 NOR2_502(n1010gat,n897gat,n455gat);
  NR2 NOR2_503(n1005gat,n894gat,n455gat);
  NR2 NOR2_504(n1182gat,n1180gat,n455gat);
  NR2 NOR2_505(n1757gat,n1773gat,n1769gat);
  NR2 NOR2_506(n1745gat,n1869gat,n1757gat);
  NR2 NOR2_507(n73gat,n67gat,n2784gat);
  NR2 NOR2_508(n70gat,n71gat,n2720gat);
  NR2 NOR2_509(n77gat,n76gat,n2784gat);
  NR2 NOR2_510(n13gat,n2720gat,n14gat);

endmodule
