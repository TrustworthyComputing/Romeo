module s38584(VDD,CK,g100,g10122,g10306,g10500,g10527,g113,g11349,g11388,
  g114,g11418,
  g11447,g115,g116,g11678,g11770,g120,g12184,g12238,g12300,g12350,g12368,g124,
  g12422,g12470,g125,g126,g127,g12832,g12833,g12919,g12923,g13039,g13049,
  g13068,g13085,g13099,g13259,g13272,g134,g135,g13865,g13881,g13895,g13906,
  g13926,g13966,g14096,g14125,g14147,g14167,g14189,g14201,g14217,g14421,g14451,
  g14518,g14597,g14635,g14662,g14673,g14694,g14705,g14738,g14749,g14779,g14828,
  g16603,g16624,g16627,g16656,g16659,g16686,g16693,g16718,g16722,g16744,g16748,
  g16775,g16874,g16924,g16955,g17291,g17316,g17320,g17400,g17404,g17423,g17519,
  g17577,g17580,g17604,g17607,g17639,g17646,g17649,g17674,g17678,g17685,g17688,
  g17711,g17715,g17722,g17739,g17743,g17760,g17764,g17778,g17787,g17813,g17819,
  g17845,g17871,g18092,g18094,g18095,g18096,g18097,g18098,g18099,g18100,g18101,
  g18881,g19334,g19357,g20049,g20557,g20652,g20654,g20763,g20899,g20901,g21176,
  g21245,g21270,g21292,g21698,g21727,g23002,g23190,g23612,g23652,g23683,g23759,
  g24151,g24161,g24162,g24163,g24164,g24165,g24166,g24167,g24168,g24169,g24170,
  g24171,g24172,g24173,g24174,g24175,g24176,g24177,g24178,g24179,g24180,g24181,
  g24182,g24183,g24184,g24185,g25114,g25167,g25219,g25259,g25582,g25583,g25584,
  g25585,g25586,g25587,g25588,g25589,g25590,g26801,g26875,g26876,g26877,g27831,
  g28030,g28041,g28042,g28753,g29210,g29211,g29212,g29213,g29214,g29215,g29216,
  g29217,g29218,g29219,g29220,g29221,g30327,g30329,g30330,g30331,g30332,g31521,
  g31656,g31665,g31793,g31860,g31861,g31862,g31863,g32185,g32429,g32454,g32975,
  g33079,g33435,g33533,g33636,g33659,g33874,g33894,g33935,g33945,g33946,g33947,
  g33948,g33949,g33950,g33959,g34201,g34221,g34232,g34233,g34234,g34235,g34236,
  g34237,g34238,g34239,g34240,g34383,g34425,g34435,g34436,g34437,g34597,g34788,
  g34839,g34913,g34915,g34917,g34919,g34921,g34923,g34925,g34927,g34956,g34972,
  g35,g36,g44,g5,g53,g54,g56,g57,g64,g6744,g6745,g6746,g6747,g6748,g6749,g6750,
  g6751,g6752,g6753,g72,g7243,g7245,g7257,g7260,g73,g7540,g7916,g7946,g8132,
  g8178,g8215,g8235,g8277,g8279,g8283,g8291,g8342,g8344,g8353,g8358,g8398,g84,
  g8403,g8416,g8475,g8719,g8783,g8784,g8785,g8786,g8787,g8788,g8789,g8839,
  g8870,g8915,g8916,g8917,g8918,g8919,g8920,g90,g9019,g9048,g91,g92,g9251,
  g9497,g9553,g9555,g9615,g9617,g9680,g9682,g9741,g9743,g9817,g99);
input VDD,CK,g35,g36,g6744,g6745,g6746,g6747,g6748,g6749,g6750,g6751,g6752,
  g6753,g84,
  g120,g5,g113,g126,g99,g53,g116,g92,g56,g91,g44,g57,g100,g54,g124,g125,g114,
  g134,g72,g115,g135,g90,g127,g64,g73;
output g7243,g7245,g7257,g7260,g7540,g7916,g7946,g8132,g8178,g8215,g8235,g8277,
  g8279,g8283,g8291,g8342,g8344,g8353,g8358,g8398,g8403,g8416,g8475,g8719,
  g8783,g8784,g8785,g8786,g8787,g8788,g8789,g8839,g8870,g8915,g8916,g8917,
  g8918,g8919,g8920,g9019,g9048,g9251,g9497,g9553,g9555,g9615,g9617,g9680,
  g9682,g9741,g9743,g9817,g10122,g10306,g10500,g10527,g11349,g11388,g11418,
  g11447,g11678,g11770,g12184,g12238,g12300,g12350,g12368,g12422,g12470,g12832,
  g12919,g12923,g13039,g13049,g13068,g13085,g13099,g13259,g13272,g13865,g13881,
  g13895,g13906,g13926,g13966,g14096,g14125,g14147,g14167,g14189,g14201,g14217,
  g14421,g14451,g14518,g14597,g14635,g14662,g14673,g14694,g14705,g14738,g14749,
  g14779,g14828,g16603,g16624,g16627,g16656,g16659,g16686,g16693,g16718,g16722,
  g16744,g16748,g16775,g16874,g16924,g16955,g17291,g17316,g17320,g17400,g17404,
  g17423,g17519,g17577,g17580,g17604,g17607,g17639,g17646,g17649,g17674,g17678,
  g17685,g17688,g17711,g17715,g17722,g17739,g17743,g17760,g17764,g17778,g17787,
  g17813,g17819,g17845,g17871,g18092,g18094,g18095,g18096,g18097,g18098,g18099,
  g18100,g18101,g18881,g19334,g19357,g20049,g20557,g20652,g20654,g20763,g20899,
  g20901,g21176,g21245,g21270,g21292,g21698,g21727,g23002,g23190,g23612,g23652,
  g23683,g23759,g24151,g25114,g25167,g25219,g25259,g25582,g25583,g25584,g25585,
  g25586,g25587,g25588,g25589,g25590,g26801,g26875,g26876,g26877,g27831,g28030,
  g28041,g28042,g28753,g29210,g29211,g29212,g29213,g29214,g29215,g29216,g29217,
  g29218,g29219,g29220,g29221,g30327,g30329,g30330,g30331,g30332,g31521,g31656,
  g31665,g31793,g31860,g31861,g31862,g31863,g32185,g32429,g32454,g32975,g33079,
  g33435,g33533,g33636,g33659,g33874,g33894,g33935,g33945,g33946,g33947,g33948,
  g33949,g33950,g33959,g34201,g34221,g34232,g34233,g34234,g34235,g34236,g34237,
  g34238,g34239,g34240,g34383,g34425,g34435,g34436,g34437,g34597,g34788,g34839,
  g34913,g34915,g34917,g34919,g34921,g34923,g34925,g34927,g34956,g34972,g24168,
  g24178,g12833,g24174,g24181,g24172,g24161,g24177,g24171,g24163,g24170,g24185,
  g24164,g24173,g24162,g24179,g24180,g24175,g24183,g24166,g24176,g24184,g24169,
  g24182,g24165,g24167;

  wire g5057,g33046,g2771,g34441,g1882,g33982,g6462,g25751,g2299,g34007,g4040,
    g24276,g2547,g30381,g559,g640,g3017,g31877,g3243,g30405,g452,g25604,g464,
    g25607,g3542,g30416,g5232,g30466,g5813,g25736,g2907,g34617,g1744,g33974,
    g5909,g30505,g1802,g33554,g3554,g30432,g6219,g33064,g807,g34881,g6031,
    g6027,g847,g24216,g976,g24232,g4172,g34733,g4372,g34882,g3512,g33026,g749,
    g31867,g3490,g25668,g6005,g24344,g4235,g4232,g1600,g33966,g1714,g33550,
    g3649,g3625,g3155,g30393,g3355,g31880,g2236,g29248,g4555,g4571,g3698,
    g24274,g6073,g31920,g1736,g33973,g1968,g30360,g4621,g34460,g5607,g30494,
    g2657,g30384,g5659,g24340,g490,g29223,g311,g26881,g6069,g31925,g772,g34252,
    g5587,g30489,g6177,g29301,g6377,g6373,g3167,g33022,g5615,g30496,g4567,
    g33043,g3057,g28062,g3457,g29263,g6287,g30533,g1500,g24256,g2563,g34015,
    g4776,g34031,g4593,g34452,g6199,g34646,g2295,g34001,g1384,g25633,g1339,
    g24259,g5180,g33049,g2844,g34609,g1024,g31869,g5591,g30490,g3598,g30427,
    g4264,g21894,g767,g33965,g5853,g34645,g3321,g3317,g2089,g33571,g4933,
    g34267,g4521,g26971,g5507,g34644,g3618,g6291,g30534,g294,g33535,g5559,
    g30498,g5794,g25728,g6144,g25743,g3813,g25684,g562,g25613,g608,g34438,
    g1205,g24244,g3909,g30439,g6259,g30541,g5905,g30519,g921,g25621,g2955,
    g34807,g203,g25599,g6088,g31924,g1099,g24235,g4878,g34036,g5204,g30476,
    g5630,g5623,g3606,g30429,g1926,g32997,g6215,g33063,g3586,g30424,g291,
    g32977,g4674,g34026,g3570,g30420,g637,g5969,g6012,g1862,g33560,g676,g29226,
    g843,g25619,g4132,g28076,g4332,g34455,g4153,g30457,g5666,g5637,g6336,
    g33625,g622,g34790,g3506,g30414,g4558,g26966,g6065,g31923,g6322,g6315,
    g3111,g25656,g117,g30390,g2837,g26935,g939,g34727,g278,g25594,g4492,g26963,
    g4864,g34034,g1036,g33541,g128,g28093,g1178,g24236,g3239,g30404,g718,
    g28051,g6195,g29303,g1135,g26917,g6137,g25741,g6395,g33624,g3380,g31882,
    g5343,g24337,g554,g34911,g496,g33963,g3853,g34627,g5134,g29282,g1422,g1418,
    g3794,g25676,g2485,g33013,g925,g32981,g48,g34993,g5555,g30483,g878,g875,
    g1798,g32994,g4076,g28070,g2941,g34806,g3905,g30453,g763,g33539,g6255,
    g30526,g4375,g26951,g4871,g34035,g4722,g34636,g590,g32978,g6692,g6668,
    g1632,g30348,g5313,g24336,g3100,g3092,g1495,g24250,g6497,g6490,g1437,
    g29236,g6154,g29298,g1579,g1576,g5567,g30499,g1752,g33976,g1917,g32996,
    g744,g30335,g3040,g31878,g4737,g34637,g4809,g25693,g6267,g30528,g3440,
    g25661,g3969,g4012,g1442,g24251,g5965,g30521,g4477,g26960,g1233,g24239,
    g4643,g34259,g5264,g30474,g6329,g6351,g2610,g33016,g5160,g34643,g5360,
    g31905,g5933,g30510,g1454,g29239,g753,g26897,g1296,g34729,g3151,g34625,
    g2980,g34800,g6727,g24353,g3530,g33029,g4742,g21903,g4104,g33615,g1532,
    g24253,g4304,g24281,g2177,g33997,g3010,g25651,g52,g34997,g4754,g34263,
    g1189,g24237,g2287,g33584,g4273,g24280,g1389,g26920,g1706,g33548,g5835,
    g29296,g1171,g30338,g4269,g21895,g2399,g33588,g3372,g31886,g4983,g34041,
    g5611,g30495,g3661,g4572,g29279,g3143,g25655,g2898,g34795,g3343,g24269,
    g3235,g30403,g4543,g33042,g3566,g30419,g4534,g34023,g4961,g28090,g6398,
    g31926,g4927,g34642,g2259,g30370,g2819,g34448,g4414,g26946,g5802,g2852,
    g34610,g417,g24209,g681,g28047,g437,g24206,g351,g26891,g5901,g30504,g2886,
    g34798,g3494,g25669,g5511,g30480,g3518,g33027,g1604,g33972,g4135,g28077,
    g5092,g25697,g4831,g28099,g4382,g26947,g6386,g24350,g479,g24210,g3965,
    g30455,g4749,g28084,g2008,g33993,g736,g802,g3933,g30444,g222,g33537,g3050,
    g25650,g5736,g31915,g1052,g25625,g58,g30328,g2122,g30366,g2465,g33593,
    g6483,g25755,g5889,g30502,g4495,g33036,g365,g25595,g4653,g34462,g3179,
    g33024,g1728,g33552,g2433,g34014,g3835,g29273,g6187,g25748,g4917,g34638,
    g1070,g30341,g822,g26899,g6023,g914,g30336,g5339,g5335,g4164,g26940,g969,
    g25622,g2807,g34447,g5424,g25709,g4054,g33613,g6191,g25749,g5077,g25704,
    g5523,g33053,g3680,g3676,g6637,g30555,g174,g25601,g1682,g33971,g355,g26892,
    g1087,g1083,g1105,g26915,g2342,g33008,g6307,g30538,g3802,g6159,g25750,
    g2255,g30369,g2815,g34446,g911,g29230,g43,g34789,g3983,g1748,g33975,g5551,
    g30497,g5742,g31917,g3558,g30418,g5499,g25721,g2960,g34622,g3901,g30438,
    g4888,g34266,g6251,g30540,g6358,g1373,g32986,g25648,g157,g33960,g2783,
    g34442,g4281,g4277,g3574,g30421,g2112,g33573,g1283,g34730,g433,g24205,
    g4297,g4294,g5983,g1459,g1399,g758,g32979,g5712,g25731,g4138,g28078,g4639,
    g34025,g6537,g25763,g5543,g30481,g1582,g3736,g31890,g5961,g30517,g6243,
    g30539,g632,g34880,g1227,g24242,g3889,g30436,g3476,g29265,g1664,g32990,
    g1246,g24245,g6128,g25739,g6629,g30553,g246,g26907,g4049,g24278,g4449,
    g26955,g2932,g24282,g4575,g29276,g4098,g31894,g4498,g33037,g528,g26894,
    g5436,g25711,g16,g34593,g3139,g25654,g102,g33962,g4584,g34451,g142,g34250,
    g5331,g5831,g29295,g239,g26905,g1216,g25629,g2848,g34792,g5805,g5798,g5022,
    g25703,g4019,g4000,g1030,g32983,g3672,g3668,g3231,g30402,g25757,g1430,
    g1426,g4452,g4446,g2241,g33999,g1564,g24262,g25729,g6148,g6140,g6649,
    g30558,g110,g34848,g884,g881,g3742,g31892,g225,g26901,g4486,g26961,g4504,
    g33039,g5873,g33059,g5037,g31899,g2319,g33007,g5495,g25720,g4185,g21891,
    g5208,g30462,g2152,g18422,g5579,g30487,g5869,g33058,g5719,g31916,g1589,
    g24261,g5752,g25730,g6279,g30531,g5917,g30506,g2975,g34804,g6167,g25747,
    g4005,g2599,g33601,g1448,g26922,g3712,g25679,g2370,g29250,g5164,g30459,
    g1333,g153,g33534,g6549,g30543,g4087,g29275,g4801,g34030,g2984,g34980,
    g3961,g30451,g5770,g25723,g962,g25627,g101,g34787,g4226,g4222,g6625,g30552,
    g51,g34996,g1018,g30337,g24254,g4045,g24277,g1467,g29237,g2461,g30378,
    g5706,g31912,g457,g25603,g2756,g33019,g5990,g33623,g471,g25608,g1256,
    g29235,g5029,g31902,g6519,g29306,g4169,g28080,g1816,g33978,g4369,g26970,
    g3436,g25660,g5787,g25726,g4578,g29278,g4459,g34253,g3831,g29272,g2514,
    g33595,g3288,g33610,g2403,g33589,g2145,g34605,g1700,g30350,g513,g25611,
    g2841,g26936,g5297,g33619,g3805,g3798,g2763,g34022,g4793,g34033,g952,
    g34726,g1263,g31870,g1950,g33985,g5138,g29283,g2307,g34003,g5109,g5101,
    g5791,g25727,g25677,g4664,g34463,g2223,g33006,g5808,g29292,g6645,g30557,
    g2016,g33989,g5759,g28098,g3873,g33033,g3632,g3654,g2315,g34005,g2811,
    g26932,g5957,g30516,g2047,g33575,g3869,g33032,g3719,g31891,g5575,g30486,
    g46,g34991,g3752,g25678,g3917,g30440,g4188,g4191,g1585,g1570,g4388,g26949,
    g6275,g30530,g6311,g30542,g4216,g4213,g1041,g25624,g2595,g30383,g2537,
    g33597,g136,g34598,g4430,g26957,g4564,g26967,g3454,g3447,g4826,g28102,
    g6239,g30524,g3770,g25671,g232,g26903,g5268,g30475,g6545,g34647,g2417,
    g30377,g1772,g33553,g4741,g21902,g5052,g31903,g5452,g25715,g1890,g33984,
    g2629,g33602,g572,g28045,g2130,g34603,g4108,g33035,g4308,g475,g24208,g990,
    g1239,g31,g34596,g3412,g28064,g45,g34990,g799,g24213,g3706,g31887,g3990,
    g33614,g5385,g31907,g5881,g33060,g1992,g30362,g3029,g31875,g3171,g33023,
    g3787,g25674,g812,g26898,g832,g25618,g5897,g30518,g4165,g28079,g6974,g3281,
    g3303,g4455,g26959,g2902,g34801,g333,g26884,g168,g25600,g2823,g26933,g3684,
    g28066,g3639,g33612,g5327,g3338,g24268,g5406,g25716,g3791,g25675,g269,
    g26906,g401,g24203,g6040,g24346,g441,g24207,g5105,g25701,g3808,g29269,g9,
    g34592,g3759,g28068,g4467,g34255,g3957,g30450,g4093,g30456,g1760,g32991,
    g6151,g24348,g160,g34249,g5445,g25713,g5373,g31909,g2279,g30371,g3498,
    g29268,g586,g29224,g869,g859,g2619,g33017,g1183,g30339,g1608,g33967,g4197,
    g4194,g5283,g5276,g1779,g33559,g2652,g29255,g5459,g2193,g30368,g2393,
    g30375,g5767,g25732,g661,g28052,g4950,g28089,g5535,g33055,g2834,g30392,
    g1361,g30343,g3419,g25657,g6235,g30523,g1146,g24233,g2625,g33018,g150,
    g32976,g1696,g30349,g6555,g33067,g26900,g3385,g31883,g3881,g33034,g6621,
    g30551,g3470,g25667,g3897,g30452,g518,g25612,g3025,g31874,g538,g34719,
    g2606,g33607,g1472,g26923,g6113,g25746,g542,g24211,g5188,g33050,g5689,
    g24341,g1116,g1056,g405,g24201,g5216,g30463,g6494,g6486,g4669,g34464,g5428,
    g25710,g996,g24243,g4531,g24335,g2860,g34611,g4743,g34262,g6593,g30546,
    g2710,g18527,g215,g25591,g4411,g1413,g30347,g4474,g10384,g5308,g6641,
    g30556,g3045,g33020,g6,g34589,g1936,g33562,g55,g35002,g504,g25610,g2587,
    g33015,g4480,g31896,g2311,g34004,g3602,g30428,g5571,g30485,g3578,g30422,
    g468,g25606,g5448,g25714,g3767,g25680,g5827,g29294,g3582,g30423,g6271,
    g30529,g4688,g34028,g5774,g25724,g2380,g33587,g5196,g30460,g5396,g31910,
    g3227,g30401,g2020,g33990,g3976,g1079,g1075,g6541,g29309,g3203,g30411,
    g1668,g33546,g4760,g28085,g262,g26904,g1840,g33556,g70,g18093,g5467,g25722,
    g460,g25605,g6209,g33062,g74,g26893,g5290,g655,g28050,g3502,g34626,g2204,
    g33583,g5256,g30472,g4608,g34454,g794,g34850,g4023,g4423,g4537,g3689,
    g24272,g5381,g31906,g5685,g5681,g703,g24214,g5421,g25718,g862,g26909,g3247,
    g30406,g2040,g33569,g4999,g25694,g4146,g34628,g4633,g34458,g1157,g24240,
    g5723,g31918,g4732,g34634,g25700,g5817,g29293,g2151,g18421,g2351,g33009,
    g2648,g33603,g6736,g24355,g4944,g34268,g4072,g25691,g344,g26890,g4443,
    g3466,g29264,g4116,g28072,g5041,g31900,g5441,g25712,g4434,g26956,g3827,
    g29271,g6500,g29304,g5673,g5654,g3133,g29261,g3333,g28063,g979,g4681,
    g34027,g298,g33961,g3774,g25672,g2667,g33604,g3396,g33025,g4210,g4207,
    g1894,g32995,g2988,g34624,g3538,g30415,g301,g33536,g341,g26888,g827,g28055,
    g24238,g6077,g31921,g2555,g33600,g5011,g28105,g199,g34721,g6523,g29307,
    g1526,g30345,g4601,g34453,g854,g32980,g1484,g29238,g4922,g34639,g5080,
    g25695,g5863,g33057,g4581,g26969,g3021,g31879,g2518,g29253,g2567,g34021,
    g568,g26895,g3263,g30413,g6613,g30549,g6044,g24347,g6444,g25758,g2965,
    g34808,g5857,g30501,g1616,g33969,g890,g34440,g5976,g3562,g30433,g21900,
    g1404,g26921,g3723,g31893,g3817,g29270,g93,g34878,g4501,g33038,g287,g31865,
    g2724,g26926,g4704,g28083,g22,g29209,g2878,g34797,g5220,g30478,g617,g34724,
    g24212,g316,g26883,g1277,g32985,g6513,g25761,g336,g26886,g2882,g34796,g933,
    g32982,g1906,g33561,g305,g26880,g8,g34591,g3368,g31884,g2799,g26931,g887,
    g4912,g34641,g4157,g34629,g2541,g33598,g2153,g33576,g550,g34720,g255,
    g26902,g1945,g29244,g5240,g30468,g1478,g26924,g3080,g25645,g3863,g33031,
    g1959,g29245,g3480,g29266,g6653,g30559,g6719,g6715,g2864,g34794,g4894,
    g28087,g5677,g3857,g30435,g499,g25609,g5413,g28095,g1002,g28057,g776,
    g34439,g28,g34595,g1236,g4646,g34260,g2476,g33012,g1657,g32989,g2375,
    g34006,g63,g34847,g358,g896,g26910,g967,g21722,g3423,g25658,g283,g28043,
    g3161,g33021,g2384,g29251,g3361,g25665,g6675,g6697,g4616,g34456,g4561,
    g26968,g2024,g33991,g3451,g3443,g2795,g26930,g613,g34599,g4527,g28082,
    g1844,g33557,g5937,g30511,g4546,g33045,g3103,g3096,g2523,g30379,g24267,
    g2643,g34020,g6109,g28100,g1489,g24249,g5390,g31908,g194,g25592,g2551,
    g30382,g5156,g29285,g3072,g25644,g1242,g47,g34992,g25662,g21896,g1955,
    g33563,g6049,g33622,g3034,g31876,g2273,g33582,g6711,g4771,g28086,g6098,
    g25744,g3147,g29262,g3347,g24270,g2269,g33581,g191,g2712,g26937,g626,
    g34849,g2729,g28060,g5357,g33618,g4991,g34038,g6019,g6000,g4709,g34032,
    g6419,g31927,g6052,g31919,g2927,g34803,g4340,g34459,g5929,g30509,g4907,
    g34640,g3298,g4035,g28069,g2946,g21899,g918,g31868,g4082,g26938,g25756,
    g2036,g30363,g577,g30334,g1620,g33970,g2831,g30391,g667,g25615,g930,g33540,
    g3937,g30445,g5782,g25725,g817,g25617,g1249,g24247,g837,g24215,g599,g33964,
    g5475,g25719,g739,g29228,g5949,g30514,g6682,g33627,g6105,g28101,g904,
    g24231,g2873,g34615,g1854,g30356,g5084,g25696,g5603,g30493,g4219,g2495,
    g33594,g2437,g34009,g2102,g30365,g2208,g33004,g2579,g34018,g4064,g25685,
    g4899,g34040,g2719,g25639,g4785,g34029,g5583,g30488,g781,g34600,g6173,
    g29300,g6369,g2917,g34802,g686,g25614,g1252,g28058,g671,g29225,g2265,
    g33580,g6283,g30532,g6365,g5320,g6459,g25760,g901,g25620,g5527,g33054,
    g4489,g26962,g1974,g33564,g1270,g32984,g4966,g34039,g6415,g31932,g6227,
    g33065,g3929,g30443,g5503,g29291,g4242,g24279,g5925,g30508,g1124,g29232,
    g4955,g34269,g5224,g30464,g2012,g33988,g6203,g30522,g5120,g25708,g2389,
    g30374,g4438,g26953,g2429,g34008,g2787,g34444,g1287,g34731,g2675,g33606,
    g66,g24334,g4836,g34265,g1199,g30340,g24257,g5547,g30482,g3782,g25673,
    g6428,g31929,g2138,g34604,g2338,g33591,g4229,g6247,g30525,g2791,g26929,
    g3949,g30448,g1291,g34602,g5945,g30513,g5244,g30469,g2759,g33608,g6741,
    g33626,g785,g34725,g1259,g30342,g3484,g29267,g209,g25593,g6609,g30548,
    g5517,g33052,g2449,g34012,g2575,g34017,g65,g34785,g2715,g24263,g936,g26912,
    g2098,g30364,g4462,g34254,g604,g34251,g6589,g30560,g1886,g33983,g6466,
    g25752,g6346,g429,g24204,g1870,g33980,g4249,g34631,g6455,g28103,g3004,
    g31873,g1825,g29243,g6133,g25740,g1008,g25623,g4392,g26950,g5002,g3546,
    g30431,g5236,g30467,g1768,g30353,g4854,g34467,g3925,g30442,g6509,g29305,
    g732,g25616,g2504,g29252,g1322,g4520,g6972,g2185,g33003,g37,g34613,g4031,
    g4027,g2070,g33570,g4812,g6093,g33061,g968,g21723,g4176,g34734,g24275,
    g4405,g4408,g872,g6181,g29302,g6381,g24349,g4765,g34264,g5563,g30484,g1395,
    g25634,g1913,g33567,g2331,g33585,g6263,g30527,g50,g34995,g3945,g30447,g347,
    g5731,g31914,g4473,g34256,g1266,g25630,g5489,g29290,g714,g29227,g2748,
    g31872,g5471,g29287,g4540,g31897,g6723,g6605,g30562,g2445,g34011,g2173,
    g33996,g4287,g21898,g2491,g33014,g4849,g34465,g2169,g33995,g2283,g30372,
    g6585,g30545,g121,g30389,g2407,g33590,g2868,g34616,g2767,g26927,g1783,
    g32992,g3310,g1312,g25631,g5212,g30477,g4245,g34632,g645,g28046,g4291,g79,
    g26896,g182,g25602,g1129,g26916,g2227,g33578,g6058,g25745,g4204,g2246,
    g33579,g1830,g30354,g3590,g30425,g392,g24200,g1592,g33544,g6505,g25764,
    g6411,g31930,g1221,g24246,g5921,g30507,g106,g26889,g146,g30333,g218,g6474,
    g25753,g1932,g32998,g1624,g32987,g5062,g25702,g5462,g29286,g2689,g34606,
    g6573,g33070,g1677,g29240,g2028,g32999,g2671,g33605,g24255,g26945,g34,
    g34877,g1848,g33558,g3089,g25647,g3731,g31889,g86,g25699,g5485,g29289,
    g2741,g30388,g2638,g29254,g4122,g28074,g4322,g34450,g5941,g30512,g2108,
    g33572,g25,g15048,g1644,g33551,g595,g33538,g2217,g33005,g1319,g24248,g2066,
    g33002,g1152,g24234,g5252,g30471,g2165,g34000,g2571,g34016,g5176,g33048,
    g391,g26911,g5005,g2711,g18528,g1211,g25628,g2827,g26934,g6423,g31928,
    g4859,g34468,g424,g24202,g1274,g33542,g85,g34717,g2803,g34445,g6451,g28104,
    g1821,g33555,g2509,g34013,g5073,g28091,g1280,g26919,g4815,g6633,g30554,
    g5124,g29281,g6303,g30537,g5069,g28092,g2994,g34732,g650,g28049,g1636,
    g33545,g3921,g30441,g2093,g29247,g6732,g24354,g1306,g25636,g5377,g31911,
    g1061,g26914,g3462,g25670,g2181,g33998,g956,g25626,g1756,g33977,g5849,
    g29297,g4112,g28071,g2685,g30387,g2197,g33577,g6116,g25737,g2421,g33592,
    g1046,g26913,g482,g28044,g4401,g26948,g6434,g31931,g1514,g30344,g329,
    g26885,g6565,g33069,g2950,g34621,g4129,g28075,g1345,g28059,g6533,g25762,
    g3274,g3085,g25646,g4727,g34633,g24352,g1536,g26925,g3941,g30446,g370,
    g25597,g5694,g24342,g1858,g30357,g446,g26908,g4932,g21905,g3219,g30399,
    g1811,g29242,g3431,g25659,g6601,g30547,g3376,g31881,g2441,g34010,g1874,
    g33986,g4349,g34257,g6581,g30544,g6597,g30561,g5008,g3610,g30430,g2890,
    g34799,g1978,g33565,g1612,g33968,g112,g34879,g2856,g34793,g6479,g25754,
    g1982,g33566,g6661,g5228,g30465,g4119,g28073,g6390,g24351,g1542,g30346,
    g4258,g21893,g4818,g5033,g31904,g4717,g34635,g1554,g25637,g3849,g29274,
    g6704,g3199,g30396,g5845,g25735,g4975,g34037,g790,g34791,g5913,g30520,
    g1902,g30358,g6163,g29299,g4125,g28081,g4821,g28096,g4939,g28088,g24241,
    g3207,g30397,g4483,g3259,g30409,g5142,g29284,g5248,g30470,g2126,g30367,
    g3694,g24273,g5481,g29288,g1964,g30359,g5097,g25698,g3215,g30398,g111,
    g34718,g4427,g26952,g7,g34590,g2779,g26928,g4200,g26954,g1720,g30351,g1367,
    g31871,g5112,g19,g34594,g4145,g26939,g2161,g33994,g376,g25596,g2361,g33586,
    g21901,g582,g31866,g2051,g33000,g1193,g26918,g5401,g33051,g3408,g28065,
    g2327,g30373,g907,g28056,g947,g34601,g1834,g30355,g3594,g30426,g2999,
    g34805,g5727,g31913,g2303,g34002,g3065,g25652,g699,g28053,g723,g29229,
    g5703,g33620,g546,g34722,g2472,g33599,g5953,g30515,g25649,g6439,g33066,
    g1740,g33979,g3550,g30417,g3845,g25683,g2116,g33574,g3195,g30410,g3913,
    g30454,g34024,g1687,g33547,g2681,g30386,g2533,g33596,g324,g26887,g2697,
    g34607,g5747,g33056,g4417,g31895,g6561,g33068,g1141,g29233,g24258,g2413,
    g30376,g1710,g33549,g6527,g29308,g6404,g25759,g3255,g30408,g1691,g29241,
    g2936,g34620,g5644,g33621,g5152,g25707,g5352,g24339,g6120,g25738,g2775,
    g34443,g2922,g34619,g1111,g29234,g5893,g30503,g1311,g21724,g3267,g6617,
    g30550,g2060,g33001,g4512,g33040,g5599,g30492,g3401,g25664,g4366,g26944,
    g94,g34614,g3129,g29260,g3329,g3325,g5170,g33047,g4456,g25692,g5821,g25733,
    g6299,g30536,g3727,g31888,g2079,g29246,g4698,g34261,g3703,g33611,g1559,
    g25638,g943,g34728,g411,g29222,g25742,g3953,g30449,g3068,g25643,g2704,
    g34608,g6035,g24345,g6082,g31922,g49,g34994,g1300,g25635,g4057,g25686,
    g5200,g30461,g4843,g34466,g5046,g31901,g2250,g29249,g319,g26882,g4549,
    g33041,g2453,g33011,g5841,g25734,g5763,g28097,g3747,g33030,g2912,g34618,
    g2357,g33010,g164,g31864,g4253,g34630,g5016,g31898,g3119,g25653,g1351,
    g25632,g1648,g32988,g4519,g33616,g5115,g29280,g3352,g33609,g6657,g30563,
    g4552,g33044,g3893,g30437,g3211,g30412,g929,g21725,g5595,g30491,g3614,
    g30434,g2894,g34612,g3125,g29259,g3821,g25681,g4141,g25687,g4570,g33617,
    g5272,g30479,g2735,g29256,g728,g28054,g6295,g30535,g5417,g28094,g2661,
    g30385,g1988,g30361,g5128,g25705,g1548,g24260,g3106,g29257,g4659,g34461,
    g4358,g34258,g1792,g32993,g2084,g33992,g3061,g28061,g3187,g30394,g4311,
    g34449,g2583,g34019,g3003,g21726,g1094,g29231,g3841,g25682,g4284,g21897,
    g3763,g28067,g3191,g30395,g4239,g21892,g3391,g31885,g4180,g691,g28048,g534,
    g34723,g5366,g25717,g385,g25598,g2004,g33987,g2527,g30380,g5456,g4420,
    g26965,g5148,g25706,g4507,g30458,g5348,g24338,g3223,g30400,g4931,g21904,
    g2970,g34623,g5698,g24343,g3416,g25666,g5260,g30473,g1521,g24252,g3522,
    g33028,g3115,g29258,g3251,g30407,g1,g26958,g4628,g34457,g1996,g33568,
    g25663,g4515,g26964,g4300,g34735,g1724,g30352,g1379,g33543,g24271,g12,
    g30326,g1878,g33981,g5619,g30500,g71,g34786,g59,g29277,I28349,g28367,
    g19408,g16066,I21294,g18274,g13297,g10831,g19635,g16349,g32394,g30601,
    I19778,g17781,g9900,g11889,g9954,g13103,g10905,g17470,g14454,g23499,g20785,
    g6895,g9797,g31804,g29385,g6837,I15824,g20066,g17433,g33804,g33250,g20231,
    g17821,I19786,g17844,g24066,g21127,g11888,g10160,g9510,I22692,g21308,
    g12884,g10392,g22494,g19801,g9245,I13031,g8925,I12910,g34248,I32243,g10289,
    g11181,g8134,I20116,g15737,g7888,g9291,g28559,g27700,g21056,g15426,I33246,
    g34970,g10288,I13718,g8224,g21611,I21210,I17932,I21285,I12530,g16521,
    g13543,I22400,g19620,g23611,g18833,g10571,g10233,g17467,g14339,g17494,
    g10308,g27015,g26869,g23988,g19277,g23924,g18997,g12217,I15070,g14571,
    I16688,g32318,g31596,g32446,g14308,I16471,I24041,g22182,I14935,g9902,
    g34778,I32976,g20511,g17929,g26672,g25275,g11931,I14749,I20816,g23432,
    g21514,I18165,g13177,I18523,g14443,g21271,I21002,I31776,g33204,g23271,
    g22155,g19074,I22539,g19606,I32231,g34123,I32988,g9259,I15190,g17782,
    I18788,I12483,g9819,I16969,g13943,g32540,g30614,g25027,I24191,g19711,
    g17062,g22170,g19210,g13190,g10939,g7297,g17419,g14965,g20660,g17873,
    g16861,I18051,g21461,g15348,g10816,I14054,g28713,g27907,g15755,g13134,
    g23461,I24237,g23823,g34945,g34933,I12779,g31833,I18006,g13638,I20035,
    g15706,I17207,g13835,g30999,g29722,g25249,g22228,g9488,g19537,g15938,
    g17155,I18205,I16855,g10473,g15563,I17140,g23031,g30090,g29134,g30998,
    g29719,g25248,g23650,g20653,g7138,g16099,g13437,g34998,g34981,g23887,
    g25552,g22594,g20916,g18008,g27084,g26673,g30182,I28419,g7963,g10374,g6903,
    I32763,g34511,g17614,g19492,g22167,g22194,I21776,g7109,g7791,I12199,g34672,
    I32800,g16777,I18003,g20550,g15864,g23529,g20558,g6854,g18930,g15789,
    g13024,g11900,g32902,g30673,g6941,g12110,I14970,g32957,g31672,g9951,g32377,
    g30984,g12922,g12297,g23528,g12321,g9637,g28678,g27800,g32739,g30735,
    g21393,g17264,g23843,g19147,g26026,I25105,g25081,g22342,g20085,g16187,
    g23393,g20739,g19750,g16326,I28594,g24076,g19984,g24085,g20857,g17589,
    g14981,g20596,I20690,g34932,g34914,g23764,g25786,g24518,I25869,g25851,
    g32738,g31376,g32562,g32645,g30825,g14669,g12301,g20054,g17328,I26337,
    g26835,g24054,g19919,I20130,g15748,g17588,g14782,g17524,g14933,I18600,
    g23869,g32699,g31528,g6989,I28576,g28431,I28585,g30217,I15987,g12381,
    g14668,g12450,g25356,g22763,g24431,g22722,g29725,g28349,I15250,g9152,
    g28294,g27295,g8945,g10489,g11987,I14833,g13625,g10971,I25161,g24920,
    g17477,g14848,g23868,g32698,g31812,g11250,g7502,g25380,g23776,I32550,
    g34398,g7957,g13250,I15811,g20269,g15844,g34505,g34409,g7049,g20773,I20830,
    g25090,g23630,g6958,g20268,g14424,g11136,I32881,g12417,g7175,g25182,g12936,
    g12601,g20655,I20753,g8340,I16231,g21225,g17428,g24156,I23312,g23259,
    g21070,g24655,g23067,I12109,I18063,g14357,g7715,g29744,g8478,g20180,g17533,
    g17616,g14309,g20670,I29447,g30729,g10830,g10087,g34134,g22305,I23384,
    g32632,g31070,g31795,I29371,g9594,g6829,g7498,g23258,g20924,g26811,g25206,
    I16590,g11966,g10544,I13906,g15573,I17154,I27492,g27511,g9806,g14544,
    I16663,I14653,g9417,I33044,g34775,I16741,g25513,g23870,g32661,g20993,
    g15615,g32547,g32895,g8876,I12855,g24839,g23436,g23244,I22343,g24993,
    g22384,g22177,g16162,g11855,I14671,g20667,g15224,g17466,g12983,g9887,
    I11746,g24667,g23112,g9934,g21069,g15277,g25505,g34433,I32470,g34387,
    g34188,g10042,g24131,g21209,g32481,g31194,I16803,I13321,g18975,g19553,
    g16782,g19862,I20233,g30097,g29118,I12884,g16629,g13990,I16150,g10430,
    g21657,g17657,g16472,g14098,I20781,g21068,g14255,I21477,g18695,I16391,
    g32551,g32572,g23375,I24781,g24264,I33146,g34903,g7162,g25212,g7268,I11740,
    g7362,g12909,g10412,g9433,g26850,I25576,g12543,g17642,g14691,g20502,g15373,
    g10678,I13990,I22725,g21250,I13740,g23879,I20647,g23970,g34343,g34089,
    g20210,g16897,I22114,g19935,g12908,g10414,g20618,g11867,I14679,g11894,
    I14702,I11685,g8310,g23878,g21337,g15758,g20443,g15171,g10383,g6978,g23337,
    g19757,g17224,g9496,g14383,I16535,g17733,g14238,I16526,g8663,g10030,g23886,
    g21468,I18614,g32490,g10093,g18884,g27242,g26183,I14576,g8791,g11714,g8107,
    g22166,g11450,I14455,I17114,g14358,I27192,g27662,g23792,g23967,g23994,
    g32784,g9891,I18320,g13605,g28037,g26365,g8002,g9337,g9913,g32956,g18215,
    g11819,g7717,g11910,g10185,g14065,g11048,g7086,g13707,g11360,g31829,g32889,
    g11202,I14267,g8236,g33920,I31786,I21254,g16540,g24039,g21256,I24759,
    g21425,g15509,I27579,I17744,g14912,g23459,I16917,g10582,g20038,g23425,
    g20751,g31828,g32888,g10108,g25097,g32824,g10219,g13055,I15682,g9807,
    I30901,g32407,g19673,g16931,g24038,g21193,g14219,g19397,g16449,g21458,
    g6849,I15590,g11988,g28155,I26664,I13762,g6755,g13070,g11984,g23458,I22583,
    g32671,I21036,g17221,g34229,g33936,g10218,I18034,g13680,g16172,g13584,
    g20601,g21010,g15634,g11986,I14830,g7470,g17476,g14665,g17485,I18408,
    I16077,I14745,g10029,g11741,g10033,g22907,g20453,g23545,g21562,g23444,
    I22561,g25369,g32931,g30937,g33682,I31515,g6900,g19634,g19872,g17015,
    g34716,I32878,I20542,g16508,I25598,g25424,g8928,g29812,g28381,I28241,
    g28709,g12841,g10357,I21934,g10981,g9815,g8064,g13017,I20913,g16964,g23086,
    g20283,I32815,g34470,g30310,g28830,g8899,g11735,g8534,g29371,I27735,I11908,
    g9692,g13877,g11350,I32601,g34319,I12767,I23351,g24791,g23850,I13166,
    I16102,g26681,g25396,g20168,g9154,I12994,g25133,g23733,I33167,I26309,
    g26825,g9354,g27014,g25888,I27564,g28166,I23348,g23322,I22425,g32546,
    g31170,g9960,g22519,g22176,I16401,g26802,I25514,g28119,g27008,g12835,
    g10352,g7635,g14277,I16455,g20666,g13018,I15636,g10520,g32024,I29582,
    g25228,g23828,I19802,g15727,g19574,g16826,g7766,I12189,g19452,g6819,I19857,
    g16640,g22154,g7087,I33297,g35000,g25011,g32860,I18891,g16676,g7487,I33103,
    g34846,g8237,g18953,g16077,I14761,g7753,g19912,I18460,g21561,g15595,I12183,
    g21656,g17700,g6923,g26765,g25309,I25680,g25641,g22935,g17092,g14011,
    g34944,g10037,I32791,g34578,g32497,g21295,g23353,g29507,g28353,I32884,
    g34690,g8844,I12826,g11402,g7594,g17518,g14918,g26549,I25391,g17154,g14348,
    g22883,g20391,g20556,g15483,I22989,g17637,g12933,g20580,g26548,g25255,
    g10419,g8821,g11866,g9883,g11917,I14727,g32700,g31579,I26687,g27880,g32659,
    g21336,g17367,g32625,g6804,g23336,I32479,g34302,g19592,g34429,I32458,
    g10155,g10418,g8818,g12041,I14905,g32658,g19780,g16739,g13223,g12430,
    I16660,g34428,I32455,I21074,g17766,g23966,g22215,g28036,g27237,g26162,
    g32943,g31710,g20110,g11706,I14579,g24084,g20720,g16738,I17956,g9761,
    g13706,g11280,g16645,g13756,g12465,g7192,I11992,g24110,g20922,I20891,
    g27983,g26725,g20321,g23017,g32644,g33648,I31482,I21238,I32840,g6870,g9828,
    g20179,g17249,g34549,I32617,g8948,g20531,g15907,I15600,I23381,g16290,
    g13260,g32969,g13280,I15846,g6825,g33755,I31610,g17501,I18434,g7369,g27142,
    g26105,g8955,g20178,g16971,g10194,g19396,g16431,I18504,g13624,g10951,
    I14241,g8356,I21941,g18918,I23378,I16371,g32968,g19731,g17093,g29920,
    g28824,g34504,g34408,g29358,I27718,g7868,I15102,I26195,g26260,I11835,g9746,
    I13326,g20373,g32855,g23289,g24685,g23139,g24373,g22908,I33024,g34783,
    g8150,g10401,g7041,g22906,I20750,I16596,g12640,g34317,g34115,g8350,g18908,
    g16100,g32870,g31021,g7535,g32527,I13007,g8038,I12360,g10119,I24474,g22546,
    g16632,g8438,g23571,g28693,g27837,g23308,g21024,g31794,I29368,g31845,g8009,
    I31497,g33187,g7261,g24417,g22171,g33845,I31694,g10118,I19775,g17780,g9932,
    g28009,I26516,g16661,I17507,g13416,g25549,g13876,g11432,g13885,g10862,
    g32503,g23495,I22622,I31659,g33219,I16829,g32867,g32894,I31625,g33197,
    g14616,I16733,g34245,I32234,I32953,g34656,g8836,g30299,g28765,g6887,g23816,
    g25548,g22550,g34323,g34105,g34299,g34080,I32654,g34378,g22139,I21722,
    I12893,g24964,I24128,g7246,g26856,I25586,g13763,g14276,I16452,I29182,
    g34582,g32581,g32714,g32450,g31591,g10053,g23985,g22138,g21370,g15739,
    g13284,I26705,g27967,I32967,g16677,g20587,g32707,g32819,g9576,g31832,
    I20982,g16300,g23954,I23099,g24587,g8229,g9716,I22788,g18940,I26679,g27773,
    g12863,g10371,g8993,g15562,g14943,g32818,g10036,g32496,g19787,g17096,
    g16127,g8822,g10177,g20909,g17955,g20543,I13684,I29441,g9848,g21669,I21230,
    I19837,g17415,g14797,g6845,I15550,g32590,g31154,g9699,g9747,I13329,g24117,
    g24000,I33197,g34930,g23260,g19743,g17125,I14584,g9766,g33926,I31796,
    g25245,g34697,g34545,g26831,g24836,g20569,I20840,g17727,I33285,g23842,
    g32741,g13314,g10893,g23384,g25299,g32384,g31666,I19831,g16533,g33388,
    g32382,I18252,I16502,g20568,g23489,g25533,I15717,g19769,g16987,g24568,
    g22942,g20242,g16308,g25298,g23760,g11721,g10074,g7689,I12159,g29927,
    g28861,I17121,g14366,g34512,g34420,g21424,g23559,g13596,g23525,g23488,
    g28675,g27779,g23016,I32909,g34712,g7216,g11431,g7618,g12952,I15572,g23558,
    g13431,I15932,g32801,g14630,g12402,g32735,g24123,g21143,g32877,g7028,
    I11785,I30686,g32381,g8895,g10166,g17576,g14953,g17585,g14974,g20772,g9644,
    g22200,g23893,I15773,g11269,g7516,I15942,g14166,g8620,g19881,g15915,g8462,
    g25232,g29491,I27777,g7247,g20639,I17173,g13716,I18101,I16468,g12760,
    g23544,g23865,I12046,g32695,I31581,g33164,g11268,g7515,g20230,I20499,
    g12790,g7097,g17609,g14817,g29755,I28002,g7564,g20638,I18509,g9818,g13655,
    g10573,g34316,g34093,g17200,I18238,g32526,g20265,g29981,g28942,g6815,
    I12787,g12873,g10380,I22028,g20204,I29211,g30298,I12776,I18872,g13745,
    I23333,g22683,g30989,g29672,g33766,I31619,g19662,g17432,g21610,I16613,
    g23610,g10570,g9021,g34989,I33267,g8249,I20562,g32457,g21189,g24992,g22417,
    I33070,g34810,g20510,g17226,g23189,g20060,g11930,g9281,I15238,g26736,
    g25349,g9186,I13010,g17745,g14978,g34988,I33264,g22973,g20330,g34924,
    I33164,g6960,g9386,I15667,g12143,I32639,g34345,I20999,g32866,g32917,g23270,
    g19482,g21678,I18813,g12834,g10349,g20579,g34432,I32467,g7308,g11965,
    I14797,g8085,I12382,g9599,g19710,g17059,g18983,g24579,g34271,g34160,g19552,
    g16856,g21460,g15628,g21686,g9274,g20578,g26843,I25567,g23460,g23939,
    g21383,g19779,I19843,g16594,g9614,I33067,g34812,I18647,g12021,g9543,g10823,
    g20586,g23030,g32706,g23938,g32597,I18574,g13075,g25316,g8854,g21267,
    g15680,g24586,I32391,g34153,g23267,g20097,g9821,I13236,g14563,g34145,
    I32096,I16168,g24842,g32689,g15824,I17324,g20442,g10382,I18912,g15050,
    I22240,g20086,g32923,g33451,g32132,g19786,g10142,I17857,g12614,g9935,
    g22761,g9280,I13054,g10519,g9326,g34736,I32904,g10176,I16479,g27320,I26004,
    I18135,g32688,g32624,g21681,g13279,I15843,I16217,I21115,g15714,g16658,
    g14157,I22604,g10518,g9311,g10154,g12905,g10408,g20615,g33246,g32212,g9083,
    g23875,g25080,g23742,g24116,I16639,g23219,I22316,I28591,g13278,g10738,
    g26709,g25435,I29969,g30991,g8219,g27565,g26645,I17491,I16486,g11204,
    g20041,g15569,g9636,g22214,g7827,g12122,g9705,g20275,g24041,g19968,g19998,
    g8431,g11468,g7624,g16644,I17842,I15663,g8812,I12805,g22207,I21787,g6828,
    g19672,g34132,g33831,I18333,I12890,g29045,g34960,I33218,g11038,g8632,
    g16969,g14262,g6830,g17013,I18350,g8005,g20237,g17213,g21160,g17508,g7196,
    I11860,g11815,g7582,g8405,I12572,g9187,g16968,I27552,g28162,I15677,g31859,
    I32116,g33937,g20035,g16430,g31825,g32876,g32885,g34161,g33851,g16197,
    g13861,g24035,g20841,g11677,g21455,I12003,g8286,g8765,I18313,g31858,g13975,
    g32854,g7780,g16527,g14048,g25198,g30259,g28463,g25529,g14215,g12198,
    g32511,g23915,g32763,I15937,g11676,I17395,I28434,g28114,g30087,g29121,
    g11143,g8032,g19961,g26810,g25220,I29894,g31771,I14033,g8912,g34471,g34423,
    g9200,g25528,g21273,g31844,I31597,g8733,g19505,g23277,I22380,g7018,g8974,
    I12930,I11726,I32237,g34130,I17633,g13258,g32660,g7418,I13726,g9003,g6953,
    g7994,I12336,g29997,g29060,g11884,g8125,g21467,I16676,g10588,g25869,g25250,
    g6956,g23494,I22619,g26337,g24818,I32806,g34585,g8796,I32684,g34430,g32456,
    g34244,I33300,g35001,g20130,I22000,g13410,I15921,g21037,g24130,g20998,
    g32480,g10083,g10348,g32916,g10887,g12891,g10399,g8324,g26792,g25439,
    g20523,I16417,I21013,g15806,g32550,I13252,g23984,g18952,g16053,I23339,
    g30068,g29157,I33020,g31227,g17683,g15027,g23419,g34068,g33728,g21352,
    g16322,g13015,g11875,g8540,g23352,I24445,g25225,g23802,g21155,g15656,
    I33109,g21418,g22882,g28608,g27670,g23418,g32721,g20006,I26466,g26870,
    I15556,g11928,g32596,g9223,g12109,I14967,g19433,g23170,g20046,g7197,g22407,
    g19455,I33106,g19387,I16762,g6848,g7397,I27449,g27737,g15969,I17416,I20846,
    g16923,g17296,g12108,I14964,g10139,I15223,I17612,I24396,g23453,g6855,
    g17414,g14627,g27492,g26598,g8287,g14119,g9416,I15800,g24437,g22654,g25244,
    g19343,g16136,I33282,I17098,g14336,g32773,g32942,I13037,g20703,I27576,
    I11635,g23589,g10415,I19238,g32655,g8399,g11110,g8728,g29911,g28780,g19369,
    g15995,g33377,I32446,g23524,g27091,g28184,g32670,g33120,I12026,I21100,
    g16284,g8898,g20600,I16117,I33149,g19368,I32222,g34118,g20781,g16877,
    I18071,g23477,g32734,g33645,I31477,g22759,g19857,g26817,g25242,g7631,
    g34918,g17584,g14773,I26693,g27930,g10664,I20929,g17663,g32839,g32930,
    g20372,g17847,g30079,g29097,g19412,g16489,I11903,g22758,g24372,g22885,
    g16695,g25171,g20175,I20433,g7301,I16747,g12729,I12503,g11373,g7566,g23864,
    g25886,g24537,g23022,g32667,g32694,g32838,I31550,g33698,I31539,I23369,
    g29147,g32965,g12840,g10356,g6818,g17759,g14864,g6867,g16526,g13898,g23749,
    g11607,I17228,g9880,g23313,g25994,g24575,I12523,g9537,g29950,g28896,g24063,
    g20014,g17758,g14861,g26656,g25495,g20516,I20609,g10554,g18905,g24137,
    g32487,g24516,g22670,g7751,g23285,g20887,g26680,g25300,g32619,g8259,g21305,
    g21053,g32502,g14609,I16724,g15979,I17420,g10200,g23305,g32557,g13334,
    g29151,g27858,g29172,g27020,I24787,g24266,g9978,g30322,g10608,g9155,g29996,
    g28962,I12811,g10115,g21466,g32618,I18662,g8088,g6975,I13124,g34159,g11762,
    g7964,I13483,I13606,g11964,g21036,I20910,g7441,g20209,g33661,g33895,I31751,
    g9982,g21177,I20957,g21560,I17456,g9234,I15587,g11985,g32469,I27368,g27881,
    I18482,g13350,g20208,g14745,g12423,g13216,g17141,I18191,I11750,I18248,
    g12938,g19379,g17327,g26631,g25467,g12862,g10370,g17652,g15033,I32770,
    I12451,g30295,I28540,g22332,I21838,g9542,g26364,I25327,g32468,g6821,I11655,
    g19050,I19759,g34680,I32820,g8951,g16689,g13923,g34144,I32093,g34823,
    I33037,g20542,I18089,I20584,g16280,g13330,g6984,g32038,g30934,g24021,
    g28241,g27064,g29318,g29029,g16688,g14045,I17814,g22406,g19506,g8114,
    g10184,g12040,I14902,I16579,I17626,g19386,g10805,I14046,I22785,g20913,
    I18778,g34336,g34112,g32815,g14184,g19603,g19742,g13117,g17135,g14297,
    g12904,g10410,g20614,g32601,I15569,g9554,g20436,I20569,g23874,I12837,
    g32677,g33127,g31950,g25322,I24497,g33176,I32834,g34472,I30537,g21693,
    g20607,g13569,g8650,I12896,g20320,g20073,I28832,g30301,I33131,g34906,
    g30017,g29085,g20274,g9213,I13020,g24073,g20530,g21665,I21226,g25158,
    I21744,g19338,g20593,I17754,g13494,g23665,g25783,I17355,g14591,g32937,
    g19429,I23345,g23320,g33385,I21849,g29044,g27742,g10761,g8411,g7411,g25561,
    g18891,g20565,g33212,I15814,g11129,g24122,I23399,g23450,g8136,g19730,
    g19428,g16090,g12183,I15033,I18233,g14639,g33354,g32329,I33210,g34943,
    g32791,g23476,g23485,I25555,g25241,g31824,g32884,g33888,g33346,g8594,
    g19765,g6756,I11623,g24034,g7074,I11801,g11772,I14623,g10400,g7002,g20641,
    g26816,g25260,g21454,I33279,g34986,g23555,I32607,g34358,g7474,I11980,
    I18245,g19690,g30309,g28959,g7992,g9490,I14563,g16511,g14130,g9166,g20153,
    g23570,I32274,g34195,g23914,g32479,g32666,g11293,g7527,g24153,I23303,
    I31469,g6904,g32363,I29891,I12112,g12872,g10379,I16057,g34308,g34088,g9056,
    g23907,g32478,g32015,I29571,g19504,g9456,g33931,I31807,I32464,g8228,g9529,
    g7863,g20136,I20399,g20635,I27742,g28819,I15929,g25017,g23699,g25272,
    I25594,g25531,I18897,g24136,g32486,g23239,g33426,g32017,g11841,g9800,
    I12997,I14395,g6841,g13394,g23567,g32556,g31554,I32797,g34581,I14899,
    g10198,g8033,g23238,g11510,g7633,g13510,I15981,g17812,I18810,g34816,I33030,
    g17010,g32580,g9698,g28441,g27629,g24759,I14633,g9340,g9964,g20164,g34985,
    I33255,g16709,g23941,g18091,I18879,g19128,g23382,g20682,I23336,g25289,
    I20954,g21185,g23519,I27730,g28752,g12047,g9591,g16307,g34954,g13014,
    g11872,g25023,g22457,g24891,g23231,I33143,g19626,g17409,g25288,g25224,
    g17487,g16721,g14072,I12793,g23518,g23154,I22264,g26488,I25366,g26424,
    I25356,g20575,I29438,g13007,g11852,g25308,g8195,g8137,g32922,g8891,g19533,
    g16261,g24474,g23620,g20711,I16193,I17675,I27549,g28161,g27051,I25779,
    g32531,I13847,g7266,I31791,g20327,g23935,g24711,g34669,g26830,g24411,
    g27592,g26715,g12051,g9595,g20537,g15345,g24109,g32740,g15885,I17374,g8807,
    g11615,g6875,g9619,g17507,g15030,I24331,g22976,g34668,I32788,g13116,g10935,
    g16773,g14021,I18148,g13526,g24108,I28162,g28803,g32186,I29720,g34392,
    g34202,g32676,g32685,I31491,g28399,g27074,g30195,g7400,g8859,g32953,g31327,
    g19737,g11720,I14589,I20529,g6811,I32150,g20606,g16655,g14151,g10882,g7601,
    I18104,g7092,I13634,g31658,I29242,I13872,g13041,g32654,g9843,g33658,g33080,
    g16180,g30016,g29049,g9989,I24448,g22923,g11430,g7617,g22541,I21911,g34559,
    g34384,g10407,g7063,g32800,g32936,g19697,g16886,I31486,g23215,g12820,
    I17699,g23501,g6874,I29965,g31189,I32109,g33631,I21033,g20381,I12519,
    g11237,I14305,g9834,g9971,I21234,g24982,g26679,g25385,g34830,g34893,I33119,
    g9686,g22359,g19495,g8255,g17473,g14841,g20091,I22366,g24091,g7183,g8481,
    I12618,I12128,g17789,g14321,g29956,I28185,g28180,g34544,I32613,g15480,
    I17125,g27708,g22358,g32762,g9598,I23366,g8097,g32964,g29980,g28935,g7779,
    g34713,I32871,g8497,g13142,g10632,g21349,g8154,g17325,I18304,g8354,g18948,
    g15800,g7023,g31855,g10206,g14441,g14584,g9321,g7423,g9670,I22547,g25195,
    g16487,I17695,g23906,g26093,g24814,g30610,I28872,g18904,g32587,g15085,
    I17008,I32982,g34749,g23284,g19445,g10725,g7846,g21304,g25525,g34042,
    g33674,g23800,g16234,g23304,g25016,g23666,I33179,g7161,I11843,g19499,
    g17121,g7361,g22682,g10114,g20192,g17268,g9253,I16821,I17661,g13329,g27929,
    I26448,g25558,g23566,g32909,g10082,g32543,g34270,I27232,g27993,g19498,
    g16752,g33875,g7051,I11793,g10107,g22173,I21757,g34124,g33819,g9909,g12929,
    g12550,g25830,g24485,g27583,g26686,g20663,g27928,g25893,g24541,I12761,
    g7451,g32908,g6982,g7327,g24522,g22689,I31748,g11165,I14222,g8112,g8218,
    g34939,g34922,g9740,g8267,g25544,g32569,I32388,g29190,g27046,g34480,I18276,
    g14744,g12578,g16286,I17615,g21139,g21653,g26837,g24869,I12120,g34938,
    g34920,g23653,g9552,g15655,g13202,I31800,g7017,g32568,g32747,I18310,g12978,
    I20369,g17690,g18062,g21138,g24483,I23688,g19432,g30065,I11820,g23138,
    I26799,g27660,g20553,g31819,g8676,I15727,I32192,g33628,g10398,g6999,I18379,
    g13012,g14398,I16555,g10141,g10652,g10804,g9772,g6800,I13152,g9687,I13287,
    g31818,g32814,g20326,g23333,g13222,g10590,g19753,g16601,I17783,I18752,
    I17879,I22889,g18926,g20536,g18065,g20040,g17271,I20412,g16213,g32751,
    g32807,g32772,I26952,g32974,g8830,g24040,g20702,g30218,g28918,g25188,
    g23909,g32639,g20904,g14562,g23963,g19650,g28033,g8592,g7072,g14332,I16492,
    I11691,g28954,g32638,g7472,g19529,I15382,g22927,I22128,g9860,g10406,g7046,
    I24228,g22409,g20564,g10361,g25296,g7443,g8703,I12709,g14406,g12249,g19528,
    g19696,I32119,g25267,g19330,g17326,I17181,I17671,I29363,g23585,g32841,
    g11236,g8357,I21291,g18273,g7116,g22649,g19063,I13875,I26430,g19365,g16249,
    g20673,g32510,g9691,g31801,I15821,I12056,I23393,g34708,g14833,g11405,
    g19869,g21609,g19960,g23609,g24397,g29339,g28274,g12881,g10388,g7565,
    g22903,g13175,g10909,I33137,I16593,g10498,I25115,g32579,g8068,I32621,
    g34335,g23312,I31569,I28301,g29042,I24393,I27271,g27998,g21608,g24062,
    g20509,g23608,I32158,g9607,g24509,g32578,g32835,g33695,g34277,g25218,
    g23949,g9962,g11790,I14630,g14004,g11149,g17648,g15024,g20508,g9158,I26296,
    g17491,g22981,g20634,I21029,g15816,g21052,g28163,I26682,g8677,g25837,
    g25064,g7533,g19709,g32586,I22211,g21463,g9506,I18555,I32693,g7697,g10613,
    g23745,g20900,I22024,g19350,g32442,g31213,I31814,g33149,g19471,g30037,
    g12890,g10397,g16580,g23813,g7596,I12070,g33228,g16223,g10273,I13708,
    g33457,I30989,I32062,g33653,g10106,I11743,g22845,I12887,g34984,I33252,
    g32615,I15834,g11164,g13209,g8848,g20213,I15208,g33917,I31779,g21184,
    g34419,g34151,g21674,g10812,I14050,g32720,g30155,I28390,I12563,g28325,
    g27463,g12779,g9444,g22898,g9174,g34418,g34150,g17794,g26836,g24866,I18835,
    g9374,g20574,g20452,I15542,g32430,g6918,g32746,g32493,g22719,g24452,I26100,
    g7936,g9985,g24047,g12778,g9856,g14676,I12764,g23732,g8241,I20793,g17694,
    g20912,g19602,g32465,g7117,I11816,I18323,g19657,g22718,g16740,g13980,
    I12132,g19068,g16031,g15169,I17094,g28121,g27093,g9284,g19375,I19863,
    g10795,g7202,I25692,g25689,g9239,g33923,g9180,g16186,g13555,I17876,g16685,
    g14038,g15733,I29936,g30606,I17658,g9380,g12945,g12467,g31624,I29218,
    g32806,g20072,g17384,g32684,g33688,I31523,g29707,g28504,g9832,I15073,
    g10109,g19878,g24051,g24072,g20982,I32675,g17718,g14776,g17521,g14727,
    g16654,g14136,g20592,I26512,I16575,g15479,g14895,g9853,I15593,g11989,g8644,
    g9020,g24756,I32452,g34241,g21400,g20780,g7922,g8119,g13530,g12641,g23400,
    g20676,g12998,g11829,g34836,I33050,g13593,g10556,g28173,g18929,g32517,
    g23013,I28572,g12233,g10338,I31586,g23214,g11122,g8751,I14301,g8571,g12182,
    I15030,g29978,g28927,g12672,g10003,g7581,g21329,g16577,g22926,g25155,
    g22472,g9559,g13565,g11006,g6971,I11737,I12808,I25005,I19704,g17653,g25266,
    g25170,g22498,g9931,g23539,g17573,g12911,g7597,g11034,g7611,g23005,g13034,
    g11920,g17247,I18259,I32051,g30022,g29001,I16606,g15580,g13242,g12932,
    g23538,g34864,g34840,g17389,g14915,g17926,I18852,I18120,g24152,I23300,
    g19458,I19927,g30313,g28843,I32921,g17612,g15014,g24396,g8211,g29067,
    I27401,g9905,g10541,g9407,g16423,g14066,g27961,g8186,g34313,g34086,I13552,
    I13857,g17324,I18301,g32523,g23009,g31854,g14541,g16216,I17557,I29909,
    g31791,I33041,g34772,g12897,g13409,I15918,g16587,I17763,g17777,g14908,
    g25194,I13779,g6868,I26584,g26943,g9630,g29150,g27886,g34276,g34058,g34285,
    I32284,g7995,g30305,g28939,I14192,g30053,g8026,g25524,I27970,g18827,g16000,
    g34053,g33683,g7479,g9300,g10359,g34474,g8426,g32475,g14359,I16515,g8170,
    g7840,g22997,g32727,g10358,g6827,g33660,I31494,g32863,g29196,g27059,I32846,
    g34502,g14535,g12318,g24405,g30036,I16512,g25119,I22819,I17425,g15740,
    g13342,I25683,g25642,g29313,g32437,I16875,g23235,g33456,I30986,g10121,
    g25118,g26693,g8280,I22816,I17118,g9973,g33916,I22111,g7356,I17819,g16747,
    g14113,g20583,g32703,I15474,g10364,g24020,g19532,g16821,g22360,g9040,
    g28648,g27693,I19671,I13672,g13474,I25882,g25776,g9969,g19783,I17111,
    g13809,g16123,g24046,I18845,g16814,g14058,g21414,g32600,g31542,g7704,
    I12167,g23515,g28604,g27759,g23882,g23414,I22525,g32781,I29204,g8106,
    g14173,g12076,I23324,g21697,g20113,g21407,g31243,g29933,I17590,g19353,
    g24113,I32929,g34649,g32952,g19144,g12811,g10319,g27971,g8187,g32821,g8387,
    g25036,g7163,g29597,g28444,g25101,g20105,g24357,g22325,g25560,I13548,g8756,
    g22220,I21802,g13303,I15869,g24105,g14331,I18031,g29689,I27954,g14029,
    g11283,g29923,g28874,g32790,g9648,g32137,g31134,g10028,g9875,g32516,g31655,
    I29233,I29579,g30565,g28262,I26785,g20640,I17801,g14936,g20769,g17472,
    g14656,I26406,g26187,I16040,g16224,I12086,g33670,I31504,I31727,g33076,
    g32873,g8046,g16510,g14008,g19364,g15825,g20768,g28633,g27687,g8514,g15079,
    g34570,I32868,g11796,g7985,g16579,g13267,g33335,I30861,I12568,I22886,
    g13174,g10741,I21766,g14330,g26941,I25689,I33134,g31839,g33839,I31686,
    I32827,g34477,g8345,g8841,I12823,g7157,g22147,g26519,I25380,g16578,I17750,
    I17148,g8763,I12749,I16564,g10429,g23435,g31667,g30142,g31838,g23082,
    g32834,g9839,g30074,g29046,g26518,g25233,g17591,I18526,g12896,g10402,
    g17776,g14905,g27011,g25917,I27561,g15568,g14984,g15747,g13307,g25009,
    I13723,g26818,I18868,g14315,I23360,g23360,g18945,g30567,g29930,I30962,
    g32021,g17147,g22858,I32690,I13149,g17754,I16847,I25677,g25008,g22432,
    g32542,I32803,g34584,I25399,g24489,g31487,I29149,g32453,I29981,g30931,
    g11192,g22151,I21734,I11620,I21162,g17292,I12144,I18709,g20662,g21399,
    g23849,g22996,g23940,g25892,g24528,g23399,g32726,g32913,g24027,g12946,
    g9618,g11663,g6905,g16615,g22844,g21163,g13522,g34941,g34926,g13663,g21398,
    g23848,g25555,g32614,g7626,g23398,g34688,g8858,g33443,I30971,g16720,g14234,
    g9282,g34675,I32809,I20650,g32607,g8016,I14119,g8757,I12746,g32905,I12580,
    g27112,g26793,g20710,g16746,g14258,g16309,g21278,I18832,g20552,g32530,
    g9693,g13483,g11270,g34978,I15862,g11215,g32593,g18932,g6985,g34884,g19687,
    I21246,g24003,g23263,I12631,g8522,g20779,g22319,I21831,g12378,g34935,
    I33189,g23332,g32565,g32464,g25239,g23972,g19954,g11949,I14773,g19374,
    g16047,g20778,g34883,g34852,g10794,g8470,I13206,g18897,I15536,g10395,g6995,
    g22227,g24778,g23286,g9804,g10262,g24081,g21406,g16684,g14223,g11948,
    g10224,I15702,g10838,g12944,g12659,g23406,g9792,g32641,g6832,I11665,g32797,
    g23962,g31815,g23361,I22464,g28032,I32482,g34304,g11702,g6928,g7778,g15579,
    I17159,g31601,I29207,g8654,g11182,g9621,g10191,g23500,g24356,g13621,g21049,
    I11896,g25185,I18151,g20380,g26083,g24809,g14191,I28883,I15564,g25092,
    g24999,g23626,g26284,g24875,I18337,g34501,g34400,g27730,g10521,I13889,
    g12857,I19348,g15084,g21048,g25154,g20090,g17058,g32635,g8880,I12861,
    g31937,g8595,I12666,g24090,g19489,g20233,I31823,g12793,g10287,I11716,
    g20182,g20651,g20672,g23004,I27495,g7475,g21221,I23390,g19559,g16129,
    g23221,I14644,g11183,g8135,g29942,g28867,g22957,I22143,g7627,g19558,I11708,
    g16523,g14041,g8612,g23613,I22748,g9518,g13191,I31607,g13062,g7526,I12013,
    g7998,g11509,g7632,g22146,g26653,g25337,g20513,g17301,g20449,g10389,g6986,
    g32891,I15872,g13933,g11419,g23947,g31479,I29139,I29248,I21006,g17120,
    g19544,g23273,g19865,I18728,g10612,I14684,g23605,g9776,g10099,g15746,
    g13121,g16475,g14107,g20448,I32309,I12954,g6983,I32651,g34375,g32575,
    g32474,g19713,g16816,g7439,g22698,I22009,g29993,g29018,g16727,g17738,
    g14813,g17645,g15018,g20505,g15588,g23812,g32711,g8130,g14701,g12351,
    I23318,g21689,g8542,I12644,g24505,g8330,g24404,g10272,I13705,g9965,g29965,
    g28903,I33034,g34769,g14251,g12308,I17916,g13087,g20026,g32537,I18078,
    g20212,g17194,g23234,g20375,g24026,g9264,I17302,I21058,g17747,g25438,g6973,
    I17314,g14078,I32449,g34127,g19679,I18086,g13856,g27245,g26209,g34653,
    g9360,g9933,g32606,g10032,I29236,g29498,g32492,g19678,I15205,g14032,g10140,
    I27546,g9050,g17427,I18364,I13802,g13574,I16024,g25073,g9780,g17366,g7952,
    g25083,g23782,g25348,g9450,I14450,g16600,I17780,g19686,g25284,I21189,
    g11912,g8989,g26576,g27774,g28147,I26654,I27558,g32750,I12016,I18125,
    g10061,I13581,g13311,I15878,g28754,I27238,g7616,I19484,g15122,g23507,
    g34845,g20433,g25566,g18896,g24149,g20387,g28370,g27528,I28866,g29730,
    I22180,g21366,g21421,g26718,g7004,I11777,g9379,g23421,g13051,g17691,g32796,
    g34894,g24097,g26608,g25334,g11592,I14537,g20104,g7647,g34664,I32782,
    I27713,g28224,g10360,g6836,g23012,g24104,g19890,g25139,I18700,I11697,g9777,
    g17481,g15005,I25541,g25180,g32840,I28597,g29374,I26880,I31474,g24971,
    g23590,I26427,g25138,g34576,g16873,g23541,g31800,g12995,g11820,g7503,g7970,
    I15906,g23473,g33800,I31642,g8056,I13317,I31820,g8456,g12880,g10387,I22131,
    I24078,g23789,I17839,g13412,g32192,g31262,g34851,I16357,I25359,g24715,
    I19799,g17817,g30312,g28970,I19813,g17952,g24368,g23788,g8155,g34312,
    g34098,g26973,g34200,g7224,g32522,g23359,I22458,g32663,g8355,I12534,g8851,
    I13057,g23321,g13009,I17131,g14384,I22502,g19376,g22980,I22153,g21434,
    g17248,I22557,g20695,g21358,g6839,g23434,g24850,I24022,g30052,I19674,
    g15932,g8964,I29913,g30605,I11626,g11413,g9100,I33155,g13413,g11737,g34052,
    g33635,g23946,g24133,g29169,I18894,g18944,g20229,g32483,g19617,g19470,
    g22181,g11691,I14570,g19915,g12831,g9569,g26732,g25389,I12030,g14510,g9541,
    g32553,g32862,I12089,g16726,I26649,g27675,g34813,I33027,g10776,g32949,
    g9332,I16709,g14785,g12629,I22286,g19446,g21682,I18224,g13793,I13276,g9153,
    I12991,g10147,g20716,g27989,g26759,I27567,g34973,I33235,g25554,I18571,
    g13074,g21291,g16620,g32536,g30184,g28144,g10355,g6816,g32948,g23291,
    g16607,g13960,g19494,g11929,g34674,I12487,g16320,g20582,g32702,g9744,g7095,
    g31000,g29737,g32757,g32904,g6988,I14866,g9748,g16530,g26400,I25351,I14742,
    g25115,I24281,g13583,I16028,g32621,g8872,g22520,I22601,g10151,g28120,
    g27108,I32228,g34122,g10172,g20627,g7892,g34934,g9558,g20379,g8057,g32564,
    I13995,g8744,g24379,g8457,I12935,g19352,I21918,g20050,I20321,g23029,g24112,
    g10367,g10394,g6994,I25028,g24484,g24050,g9901,g34692,g20189,I21784,g19638,
    g23506,g23028,I28480,g28652,g31814,g32673,g32847,g20386,I21297,g18597,
    g8971,I12927,g22860,g20000,g24386,g20603,g9511,g27736,I26356,g7738,I12176,
    g31807,g8686,g13302,g20096,g24603,g23108,g33772,I31622,g7991,I23354,g24096,
    g29922,g28837,g34142,g7244,g12887,g10420,I17143,g14412,g22497,g19513,
    g25184,g32509,g31639,I29225,g17088,I18160,g32933,I28588,g9492,I21181,
    g17413,g7340,g20681,g9600,I23671,g23202,g32508,g9574,g31638,g9864,I13424,
    g32634,g32851,g32872,g33638,g7907,g11640,I14550,g11769,g8626,g34539,g34354,
    g9714,g12843,g17497,g14879,g22987,g34328,g34096,g10059,g23927,I18842,
    g24429,g19524,g15695,g31578,g7517,g22658,I21969,g29953,g28907,g10540,g9392,
    g10058,g31841,g24428,g33641,g33391,g19477,g12869,g10376,g16164,g23649,
    g26683,g25514,g7876,I24839,g15614,g14914,g22339,g20765,g17748,g8938,I19235,
    g15078,I20495,g16283,g29800,g28363,g10203,g12868,g10377,I21480,g14203,
    g20549,g23648,I16181,I16090,g22338,g23491,g23903,g34974,I32681,g10044,
    g27709,g21604,I22580,I16651,g10542,g20548,g8519,g8740,I12735,I29199,g25013,
    g23599,g31835,g32574,I20985,g24548,I31564,I18280,g25214,I26334,I12418,
    g17644,g15002,g20504,g30100,g29131,g23563,g6940,g32912,g8606,I18865,g14314,
    g16228,g19748,g10120,g22197,g14377,g12201,I11753,g22855,g19276,g9889,
    g13027,I15647,g7110,I14660,g33442,g22870,g22527,g19546,I21860,g34683,
    g28127,g27102,g25538,g11249,I28838,g29372,g13249,g12036,g14645,I16755,
    g32383,g20129,g16606,g14110,g17197,g18880,g23767,g23794,g21395,g24129,
    g32592,g20057,g32756,g23395,g24057,g20128,g14290,I16460,g17870,g17411,
    g17527,g14741,g23899,g13003,I15609,g24128,I14271,g10072,g7824,I28925,g6996,
    g23651,g11779,g9602,I18270,g16750,g22867,I33273,g7236,g9285,g20626,I26381,
    g23898,g9500,g20323,I21250,g29117,g24626,g33430,g32421,g23191,I22289,
    g20533,g10427,g12955,I15577,g32820,g8341,g10366,g24533,g22876,g25100,
    g12879,g10381,g22714,g11786,g7549,g17503,g14892,g9184,g23521,g28181,I26700,
    g25771,I24920,g20775,g18831,g23232,g32846,g9339,g17767,g19733,I24558,
    g23777,g12878,g10386,g26758,I27749,g28917,g12337,g32731,g31806,g22202,
    g33806,I31650,g9024,g11826,I14650,g17714,g14930,g12886,g10393,g22979,
    g20737,g22496,g19510,g10403,g7040,g23440,g13999,g7222,I26479,g27994,g33142,
    g32072,g19630,g9809,g20232,g9581,g29814,I28062,I18825,g17707,g14758,I33047,
    g34776,g30206,g28436,g7928,g26744,g25400,g12967,g23861,g23573,g20248,
    g32691,g18989,g8879,I12858,g8607,g11233,g9664,I18875,g13782,g21247,g23247,
    g7064,g17818,I18822,g9672,g20697,g14226,g11618,g9077,g17496,g14683,I19345,
    g15083,g22986,g8659,g25882,g25026,g23926,I12541,g18988,I32775,g9477,g8506,
    I30766,g9523,g24995,g34759,I32935,g7785,g16522,g13889,I22745,g10572,I25534,
    g25448,I17964,g23388,g17590,g19476,g6799,g26804,g20512,I32476,I22918,
    g23534,I22665,I26451,g26862,g13932,g11534,g32929,g8587,I14839,g9689,g23272,
    g11513,g7948,g19454,g7563,g17741,g12972,g12918,I15533,I15448,g10877,g32583,
    g32928,g19570,g19712,g6997,g22150,g21280,g11897,I14705,g20277,g10490,g9551,
    g9742,g9104,I12987,g23462,I22589,g9099,I32352,g9499,g11404,g15750,g13291,
    g34940,g13505,g18887,g20445,g33323,I12064,g23032,g10385,I13805,g12598,
    g14376,g12126,g14385,I16541,I19772,g17735,g14807,g10869,g20499,g7394,
    g10980,g9051,g11026,g8434,g27013,g12086,g9654,g32787,g13026,g11018,I14619,
    g10354,I23315,g21685,I33152,g34900,g19567,g14095,g11326,g29014,g22526,
    I17569,g14564,g9754,g21061,g28126,g27122,g20498,g6802,g8284,g23061,g8239,
    g28250,g10181,I24278,g7557,g8180,I17747,g13298,g12322,I15162,g27977,g32743,
    g32827,g25082,g8591,g24056,g9613,g12901,g10404,g20611,g17526,I18469,g12977,
    g20080,g7471,g9044,I20895,g19519,g16795,g24080,g19675,g9269,g22866,g32640,
    g20432,g32769,I22461,g29116,g19518,g16239,g8507,g9983,g12656,I15620,g12038,
    I17772,g14888,g25849,g24491,g9862,I27555,g28142,g23447,g32768,g32803,
    g25399,g12295,g7139,g23362,g10190,g29041,I27385,g13620,g12823,g9206,I17639,
    I27570,g11128,I21067,g16509,g13873,I32056,g11811,g9724,I12712,g20145,
    g34833,g34049,g33678,g31821,g32881,g34755,g24031,g34781,I17704,I24455,
    g26605,g25293,g20650,g23629,g21451,g16872,I18060,I12907,I22124,g13806,
    g23472,g21062,I17128,g9534,g9729,g9961,g7438,g25263,g29983,g28977,g20529,
    g22300,I21815,g26812,I21019,g27017,g25895,g15862,g8515,g8630,g21246,g23246,
    g20528,g20696,g25135,g9927,g32662,g8300,g32027,I29585,I32461,g19577,I18667,
    g9014,g20764,I20819,g10497,g10102,I25591,g32890,g34987,I27941,g9414,g7212,
    g19439,g9660,g9946,g20132,g24365,g20869,g11963,g34947,g24132,g32482,g24960,
    g23716,g19438,g17157,g9903,g13133,g11330,g32710,I12092,g14700,g12512,
    g21355,g32552,g31834,g23355,g10658,I13979,g16323,g23859,g16311,g13273,
    g32779,I17442,g18878,I23327,g29130,I32696,g34434,I32843,g34499,g7993,
    I12333,g20709,g11011,g10274,g22854,g34951,I33232,g23858,g13011,I15623,
    g32778,g18886,I31803,g9036,g25221,I22275,g20127,g8440,g20708,I22046,g9679,
    g23172,g13251,g20087,g32786,g33726,I32960,g8123,g19566,g14338,g24087,
    I18285,g28590,g27724,g23844,g32647,g23394,I22499,g34579,g9831,g32945,
    g33436,g22660,g19140,I17136,I19012,g15060,g17763,g15011,g8666,g10060,
    I18900,g16767,g27976,g26703,g27985,g26131,I32161,g33791,g32826,g25273,
    g23978,g29863,g28410,g24043,g10197,I21300,g18598,g22456,g12976,I17188,
    g14197,g12160,g32090,g31003,g9805,g9916,g19653,I32225,g34121,I13892,I12577,
    g10411,g23420,g9749,I18177,I18560,g32651,g32672,I19789,g17793,g24069,
    I21922,g34767,g26788,g26724,g25341,g20657,g20774,g26859,g8655,g23446,
    I28908,g19636,g23227,g30012,g19415,g24068,g24375,g21059,I33249,g34971,
    g7462,g23059,g31797,g6838,g13096,g32932,g33797,g33306,g19852,g22721,g10503,
    I16626,g21058,g6809,g32513,I20864,g16960,g23058,g32449,I29977,g14503,
    g12256,g16691,g14160,g19963,g12842,g34473,g34426,I12083,g17085,I23357,
    g32897,g32961,g23203,I12819,I32997,g7788,g11429,g17721,g12915,I27738,
    g10581,I16775,g13857,I16163,g32505,g31566,g20994,g9095,g32404,I14800,
    g33136,g32057,g9037,g14714,g24994,g30325,I32994,g11793,g11428,g7615,g26682,
    g9653,g17431,I18376,I16120,g22341,g32717,g34325,g34092,I15765,I18009,
    g21281,g18977,I32970,g22156,g27830,g8172,g8278,I32473,g23902,g23301,I32364,
    I27314,g23377,g22180,g24425,g19554,g10111,g12830,g9995,g12893,g10391,
    g16583,g14069,g7392,g20919,g15756,g13315,I25146,g24911,g34946,I25562,
    g19609,g16264,I12463,g8343,I18476,g14031,g10230,g19200,I21199,g9752,g12865,
    g10372,g20010,g8282,g20918,g23645,g20875,g8566,g24010,g9917,I13473,g34648,
    g34739,g18696,g7854,g13504,g11303,g25541,g20545,g20079,g20444,g21290,
    g32723,I31672,I12415,g23290,I33182,g34910,I13374,g8334,g24079,g18562,
    I16538,g22667,g21156,g34682,I32824,I27543,g20599,g6926,g23698,g11317,
    I14346,g20078,g16846,g32433,I29961,g19745,g24078,g6754,I11617,g12705,
    g20598,g32620,I28579,g29474,I20355,g19799,g25325,g34243,g24477,g8804,
    g10150,g24086,g16743,g13986,g21427,g15731,g13326,g9364,I14079,g23427,
    I22542,g25535,g32811,I12963,g14150,g32646,g8792,I12790,g7219,g19798,I28014,
    g28158,g7640,g13144,g10019,g28157,I26670,I15626,g22210,I21792,g20322,
    g32971,g7431,I32079,g7252,I17834,g29913,g28840,g34760,I32938,g7812,I12214,
    g16769,g20159,g25121,I20867,g13626,g11273,g20532,I18414,g24159,I23321,
    g13323,g24125,I18382,g21661,I21222,g17502,g14697,g16768,g17408,g20158,
    g8113,I16498,g23403,I22512,g23547,g23895,g24158,g33750,I18092,g7405,g19732,
    g20100,I30980,I24008,g29905,g28783,g20561,g20656,I13202,I18518,I18154,
    g23226,g7765,g20680,g26648,g20144,g23715,g23481,g32850,g31796,g19761,
    I12608,g12875,I15494,g19268,g6961,I11734,g8567,I21930,g21297,I33173,g7733,
    I22422,I15697,I17873,g15017,g31840,g12218,g32896,g12837,g23127,g6927,
    g19263,g25134,g10001,g22975,I16160,I23694,g23252,g9888,g10077,g13995,
    g11261,g8593,g29153,g27937,g24966,g7073,I12799,g20631,g17815,g10597,g23490,
    g25506,g9429,g29505,g32716,g7473,g18976,I16713,g19539,g6946,I11721,g24017,
    g11512,g7634,I32752,g24364,g17677,g14882,g34491,g19773,g16482,g13464,
    g14977,g31522,I29185,g32582,g7980,I21042,g18954,g23376,g23385,I22488,
    I25095,g25265,g19538,g7069,g26990,g23889,g23354,g22169,g27956,g34770,
    I32956,I15284,g8160,g22884,g23888,g23824,I15831,g10416,g32627,g28307,
    g27306,g32959,g32925,g21181,g22168,g10157,I29444,g32958,I15316,I19719,
    g8450,g24023,g25168,g34208,g17791,g14950,g20571,g9684,g11316,g8967,g9745,
    g12075,I17436,I26925,g9639,I18906,g16963,g9338,g24571,g10231,I18083,g9963,
    g26820,g33326,g17410,g11498,I14475,I32947,g14231,g12246,g26832,g34773,
    g32603,g6831,g21222,g23931,g32742,g9309,I23306,g21673,g30990,g29676,g14790,
    g19771,g25240,g32944,I27758,I33270,I25190,g25423,g17479,g14855,g21426,
    g8179,g12037,I14893,g20495,g23426,g25903,g27984,g26737,g33702,I31545,g9808,
    g19683,I14836,g17478,g14996,g28156,I26667,I18143,g32681,g34210,g16182,
    g13846,g16651,g14005,g23520,g27155,g9759,g18830,g12367,g17486,I18411,g7898,
    g25563,g32802,g32857,g22223,g13271,g24985,g23586,g34521,g32730,g23546,
    I24215,g32793,I18653,g20374,g23211,I30644,g19882,g19414,g26701,g11753,
    I12538,g26777,g20643,g15962,I18138,g9049,g23088,g31847,g32765,g19407,
    g16268,g9449,I17679,g11031,g8609,g22922,g23860,I15650,g32690,g9575,g32549,
    I15736,g22179,I29717,g25262,g11736,g8165,g20669,I26503,g34573,I32645,g7344,
    g25899,g24997,g13736,g11313,g32548,I32687,g34431,g34247,I32240,g34699,
    I32985,g22178,g9498,g6873,g20668,I33170,g32504,g31851,g34510,g9833,I13715,
    g7259,g21659,g34777,I16476,g16717,g13951,g17531,g12836,g10351,g20195,
    I26581,g26942,g8997,g23987,g10085,g8541,g23250,I23363,g14307,I27235,g17178,
    I18214,g6869,I32973,g12477,I15295,g20525,g11234,g18939,I12411,g28443,
    I26936,g34272,g24525,g24424,g13132,g17676,g12941,g13869,g8680,g22936,
    I13623,I21486,g18727,g17953,I18861,I22327,g19367,g23339,g18938,g23943,
    I18885,g29384,g14431,g12208,I29013,g11868,g9185,g12864,g10373,g13868,
    g11493,g6917,g23338,g24893,I24060,g12749,g19435,g9162,I12950,g17417,g14804,
    I18609,g7886,g20544,g23969,g32626,g28039,I32195,I13352,g11709,g30997,
    g29702,g10156,g20713,g21060,I33291,g23060,g19908,g23968,g18875,g32533,
    g8558,g28038,I32525,g33912,I31770,g19744,I17808,g7314,g10180,I14006,I17108,
    g10175,g11471,g19345,g25099,g22369,g12012,g32775,g25388,g25324,g12900,
    g19399,g20610,g7870,g21411,g17762,g13000,g20705,g34766,g34703,g21293,
    I16010,g11148,g23411,g20734,g23527,g28187,I26710,g21335,g25534,g25098,
    g10335,g7650,g27101,g26770,g29862,g28406,g24042,g33072,g31945,I20447,
    g19398,g20679,g30321,I18360,I18131,g11043,g8561,g9086,g32737,g17216,g20270,
    g9728,g19652,g22543,g17587,g9730,g24124,g8092,I16795,g29948,g28853,g8492,
    g23503,g23894,g32697,I25786,I18674,g13101,g25032,g23639,g20383,g32856,
    I28913,g11810,g25140,g9070,g8714,g31820,g10487,g32880,g25997,g7972,g24030,
    g20267,g24093,g10502,g26776,g25498,g23714,I22571,I29228,g30314,g32512,
    g7806,g20065,g31846,g7943,g24065,g11878,I14690,g19361,g16539,I12758,g23819,
    g12874,g26754,g25766,g24439,g28479,g27654,I32678,I22302,g23257,g27009,
    g25911,g21055,g23496,g7322,g20219,g23055,g6990,g17242,g34246,g10278,g33413,
    g31971,g29847,g28395,g30591,g23111,g12009,I14862,I20937,g6888,I11701,
    g22974,g32831,g33691,I31528,g32445,I29973,g34663,g16716,g13948,g9678,
    g10039,g32499,g23986,I28851,g18984,g8623,I11809,g12892,g16582,g13915,
    g17772,g11425,g10038,g32498,I22485,I12141,g34147,g33823,I13280,g15811,
    g13125,g16310,g7096,g10815,g13458,g24160,g9305,g7496,g33929,g17638,g14838,
    g22841,g34950,g12914,g12235,g13010,g32611,g7845,g34957,g25451,g32722,
    g32924,g33928,g19947,g7195,g12907,g20617,g17416,g14956,g7395,g7891,g8651,
    g16958,g13545,g23877,g19273,g20915,I20882,g7913,I25790,g28321,g27317,
    I32837,g34498,g30996,g29694,g25246,I32106,I12135,g10143,I33288,g23019,
    g19866,I33261,g34977,g8285,I12497,g12074,I14932,I25695,g25690,g9226,I17787,
    g16742,g13983,g23196,g34844,g34737,I22564,g16096,g23018,g32753,g32461,
    I21242,g10169,g24075,g17579,g14959,g19371,g20595,g15877,g23526,g6808,
    g20494,g14169,g8139,I16289,g12107,g34242,g29912,g28827,g29311,g28998,
    g20623,I12049,g9373,g17014,g27092,g9091,g20037,g31827,g32736,g34333,g13322,
    g10918,g32887,g24623,g23076,g33827,g9491,g9822,g24037,g34152,g16429,g20782,
    g15853,g21457,g13901,g11480,g23402,g32529,g23457,g25370,g8795,g10363,
    I24400,g10217,I14593,g30318,g14363,I16521,g9283,g16428,I17668,g9369,g32528,
    g32696,g9007,g32843,g6957,g24419,g32393,g30922,I11892,g34059,g8672,g9920,
    I15144,g31803,g32764,g24155,I23309,g24418,g20266,g8477,g34540,g11823,
    I14647,g17615,g12883,g10390,g22493,g23001,g32869,I18882,g32960,g7497,
    g19421,g17720,g15045,I33056,g25688,g9582,g11336,g7620,g7960,g32868,g8205,
    g34571,g10223,g23256,I12106,I12605,g17430,I18373,g17746,g14825,g20853,
    g34044,g33675,g23923,I14409,g8364,g29152,g29846,g28391,g34169,I29002,
    g29675,g21300,I21047,g20167,g20194,g20589,g32709,g23300,g17465,g8742,
    I16246,g10084,g9415,g19541,I28548,g10110,g11631,g19473,I18909,g11017,
    g20588,g20524,g32708,I32170,I12033,I15633,I28174,I29245,g32471,g19789,
    g24524,I17488,g25227,g10874,g10531,g17684,g15036,g27438,I26130,g14179,
    g25025,g7267,I23680,g10178,g26632,g25473,g24119,g27349,g26352,g23066,
    g29185,g9721,I32855,g19434,g16626,g14133,g8273,g10685,I16489,I17653,g24118,
    g14186,g11346,g24022,g34698,g34550,g7293,g12906,g10413,I17733,g20616,
    I18114,g14509,g23876,I18758,g13023,g18874,g25044,g23675,I19661,g29929,
    g28914,I17999,I18107,g10417,I25511,g32602,g32810,I13637,g17619,g32657,
    g32774,g33778,g7828,g32955,g21511,g29928,g28871,g20704,g23511,I22640,
    g34427,g32879,g8572,I12654,g20053,g32970,g10334,g19682,g24053,g25120,
    g17523,g14732,g8712,g7592,I16544,I18849,g32878,g21660,g24466,g10762,g25562,
    g18892,g20036,g31826,g32886,I33161,I18398,g20101,g24036,g20560,I18048,
    g21456,g27585,I14827,g17475,g24101,I23684,g23230,g32792,g23456,g13976,
    g11130,I23375,g24560,I15954,g32967,g10216,g14423,I16610,g9671,g20642,
    g23480,g27415,g26382,g23916,g9030,g19760,I32305,g34209,I14381,g16512,
    g14015,I16679,g12039,g23550,g26784,g9247,I33258,g34976,g34586,g18907,
    g32459,g20064,g7953,g30572,g29945,g24064,g28579,g27714,g9564,g23307,g32919,
    g23085,g19957,g32458,g24229,g14543,g33932,I31810,g9826,g10117,g10000,
    g26824,g20874,g21054,g32918,g23243,g20630,g11842,g21431,g8903,g23431,
    g32545,g9910,g17600,g14659,g34490,I32547,g20166,g20009,g27576,g26081,
    g20665,g25547,g32599,I20744,g9638,g21269,g15506,I23342,g24665,g7716,g7149,
    g34784,g7349,g30297,g28758,g27554,g26625,g20008,I33214,I18858,g32598,
    g13016,g23942,g16205,g23341,g21268,g29194,g25226,g22137,I18829,I12437,
    g6801,g28615,g27817,g25481,I15893,I31878,g33696,g19649,I32874,g21180,
    I14663,g21670,I18221,I17938,g20555,g32817,g29317,g30072,g19491,g34181,
    g33913,g34671,g20570,g20712,g11865,g10124,g20914,g18883,g32532,g32901,
    I13694,g23335,I32665,g34386,g19755,g12921,g12228,g23839,g23930,g23993,
    g32783,g19770,g30237,g8805,g21694,g23838,g9861,g10318,I15705,g14044,g32561,
    g32656,g23965,I31459,g20239,g17128,g11705,g24074,I22769,g21277,g26860,
    I14326,g11042,g8691,g20567,g20594,g32680,g11845,g32823,g20238,g25297,
    g23746,g13255,g9827,g13189,g22542,g13679,g31811,g23487,I16629,g31646,g9333,
    g19794,I15036,g16529,g14055,g29081,g12805,g13188,g19395,g23502,I27927,
    g20382,I16201,I23372,g26700,g25429,g7258,I33079,g34809,g11686,I14567,
    g16528,g14154,g7577,g7867,g13460,g15831,g13385,g26987,g11383,g9061,g10014,
    g23443,g10073,I18795,g21279,g23279,g32966,g19633,I12172,g30088,g29094,
    g24092,I32074,I11688,g11030,g8292,g20154,g22905,g32631,g19719,g11294,g7598,
    g24154,I32594,g34298,g8037,g23278,g29999,g28973,g32364,g6767,g22593,I13360,
    g20637,g8102,g13065,g10476,g19718,g21286,g8302,g14442,g29998,g28966,I18297,
    g21306,g15582,g31850,g8579,g23306,g30311,I31817,g7975,g33850,I31701,g17530,
    g14947,g10116,g9662,g9018,I14687,I12719,I25743,g7026,g9467,g19440,I17919,
    g17122,g34126,I32067,g34659,I12770,g12013,g23815,g25640,I15837,I33158,
    g34897,g7170,g19861,g10275,g19573,g16708,g22153,g21677,g14275,g12358,
    g25546,g32571,I31561,I17249,g25211,g34657,g19389,g17532,g17641,g14845,
    g20501,I25606,g30296,g28889,g20577,g34339,g34077,g9816,I20951,g25024,
    g33716,g19612,g34296,I32297,g7280,g29897,I28128,g7939,g22136,g29961,g28892,
    g8442,g22408,g19483,g22635,g14237,g11666,g23937,g10035,g32495,g29186,
    g19777,I18344,I12899,g7544,g8164,g9381,I15617,g6976,g13138,g32816,I15915,
    g24438,g11470,g7625,g17136,I18341,g34060,g33704,g7636,g9685,I26676,g9197,
    g32687,g9397,g16602,g14101,g21410,g34197,g33812,g28231,g16774,g14024,
    g23410,g8770,I29337,g30286,g34855,g32752,g8296,I24434,g27100,g32954,g8725,
    g24083,g33378,I30904,g21666,g23479,g27599,g32643,g23363,I22470,g7187,g7387,
    g20622,g11467,g7623,g13595,g20566,g7461,g23478,g23015,g8553,g26834,I19707,
    g10130,g16171,g33944,I31829,g19061,I19762,I25530,I27573,g32669,I15782,
    g23486,g26055,g13037,g10362,g6850,g29149,g7027,I19818,g19766,g21556,g15669,
    g10165,g17575,g14921,g28137,I26638,g16967,I22331,g19417,g32668,g32842,
    I18694,I20747,g27991,g25852,g31802,g9631,g25060,g23708,g32489,g8389,I27388,
    g27698,g31857,g7446,g18200,g29811,g28376,g23223,g7514,g19360,I14424,g34714,
    g8990,g12882,g9257,g22492,g19614,g25197,g23958,g29343,g28174,g7003,I13539,
    g22303,g29043,g32559,g34315,g34085,g10475,g24138,g32525,g32488,g11170,
    g8476,g30928,g8171,g10727,I14016,g7345,g7841,g20636,I19384,I12773,g32558,
    g23084,g24636,g23121,g6826,g10222,g7191,g30055,g17606,g14999,g20852,g32830,
    g23922,g32893,I18028,g21179,g29368,g9751,g34070,g33725,g8281,g32544,g19629,
    g32865,g19451,g21178,g19472,g24963,g20664,g32713,g7536,g9585,g8297,g10347,
    I13759,g12026,g28726,g23953,g30067,g11401,g7593,g22840,g21654,g7858,g32610,
    g20576,g20585,g23654,I12061,g32705,g34094,g13477,g8745,I26929,g8138,g8639,
    g24585,g23063,I22149,g19071,g15591,I23711,g23192,g20554,g23417,g32679,
    I17650,g23936,g22647,g25202,g23932,g19776,g19785,I32103,I32963,g34650,
    g16159,g22192,g20609,I17723,g12082,g9645,g17390,g14755,g28593,g27727,
    g32678,g13022,g7522,g23334,g25055,g30019,g7115,g8808,g19754,g7315,g16158,
    g20608,g25111,g9669,g19355,g16027,g25070,g32460,g32686,g24115,g32939,
    I18903,g30018,g28987,g19950,g14063,g19370,I19917,g18088,I17852,g27965,
    g20921,g12345,g7158,g20052,g23964,g32938,g28034,I31361,g29310,g28991,
    g16680,g24052,I17104,g12940,g11744,g17522,g14927,g21423,g12399,g23423,
    g20871,g8201,g9890,g13305,g14873,I16898,g23216,I14708,g19996,g29379,g29925,
    g28820,I16135,g8449,g12804,g9011,I19851,g19394,g6846,g8575,g13036,g32875,
    g30917,I28897,g11560,g14209,g11415,g7880,g8715,g20674,g7595,I12067,g23543,
    g6803,g16966,g14291,g7537,I23396,g16631,g14208,g11563,I18262,g29944,g28911,
    g22904,g23000,I26578,g23908,I18307,g32837,g31856,g8833,g30077,g29057,g9992,
    g20732,g23569,g25196,g13064,g24732,g23042,g14453,I30992,I32699,g23568,
    g34975,g34929,g8584,g8539,g23242,g31783,g34689,g34982,g9863,I12355,g16289,
    g9480,g21123,g9713,g10607,g22847,g23814,g10320,g32617,g28575,g27711,g32470,
    g7328,g32915,g29765,g10530,g8922,g7542,g28711,I17636,g13665,g11306,g27004,
    g30102,g8362,I13744,g31831,g32201,g31509,g24013,g34768,I12151,g17183,
    g17673,g14723,I18839,g13008,I17198,I21483,g18726,g20329,g34979,g8052,
    g20207,g20539,g25001,g20005,g13485,g20328,g15867,g32595,g32467,g32494,
    g19902,g24005,I23149,g17509,I18446,g14034,g20538,g9688,g28606,g27762,g6847,
    g12692,g18882,g32623,g18991,g19739,g9976,I18443,I27677,g10153,g23841,
    I22096,g23992,g32782,g23391,g20645,g19146,g15574,g19738,g15992,g21510,
    g15647,g23510,g10409,I17976,g34955,I25579,g16954,g29129,g22213,g19699,
    g8504,g10136,g16643,g9000,g32822,g29128,I12227,g13239,g19698,g12951,g25157,
    g23578,g8070,g13594,g11012,I16438,g23014,g25537,g7512,g34660,I30983,g9760,
    g20771,g22311,g18935,g24100,g26054,g24804,g7490,g9071,g25231,g7166,g20235,
    g19427,g16292,g26510,g11941,g19366,g32853,g24683,g33736,g11519,I14999,
    g16195,I32535,g34916,I33140,g13675,I20861,g32589,g7456,I17101,g7148,g6817,
    g7649,g22592,g22756,g16525,g15571,g13211,g9924,g10474,g32588,g32524,g9220,
    g31843,g32836,I31535,g30076,g30085,g29082,g7851,I33075,g34843,g9779,g26655,
    g25492,g13637,g20515,g34307,g34087,g23041,I20388,g17724,g32477,g21275,
    g24515,g33283,g24991,g30054,g21430,g15608,g27163,g8406,g17756,g14858,
    g28140,g23430,g20902,g23493,g8635,g24407,g29697,g28336,g9977,g19481,g29995,
    g28955,g32118,g31008,g8766,g8087,I31782,g32864,g23237,I19734,g17725,g10606,
    g21340,g32749,g32616,g23340,g23983,g23684,g25480,g34942,g34928,g32748,
    g8748,g19127,g9451,g28326,g27414,I32991,I14505,g13215,g34156,g33907,g13729,
    g25550,g20441,g20584,g32704,g17429,g28040,g33708,I31555,g34890,g19490,
    g25287,g34670,I32794,I29939,g9999,g23517,g33258,g32296,g32809,g32900,
    g25307,g32466,g7118,g7619,g16124,I19487,g15125,g19385,g14582,g9103,g32808,
    g27972,g23003,g19980,g25243,I33053,g20114,I20385,I17892,I14365,g15842,
    g13469,g32560,g20435,g8373,g24114,g8091,g6772,I11629,I27784,g24082,g16030,
    g13570,g7393,g6987,g21362,g24107,g32642,g9732,I22467,g34131,g29056,g22928,
    g9753,g23523,g31810,I12493,g25773,g24453,I27481,g31657,I29239,g7971,g13304,
    g16244,I28582,g30116,I18370,g24744,g29080,g7686,g33375,g8407,I18855,g9072,
    g25156,g30304,g8059,g32733,g14192,g11385,g9472,g19931,g6856,I11682,g15830,
    g13432,g17583,g14968,g8718,I32173,g32874,g29987,g9443,g28508,I26989,g32630,
    g7121,g23863,g32693,I31616,g7670,g23222,I18367,g29342,g28188,g9316,g25930,
    g32665,g19520,g6992,g9434,g7232,g10553,g25838,g29013,I33276,g18947,g30039,
    g30306,g28796,g25131,g15705,g13217,g17302,g32892,g23347,I22444,g24135,
    g32476,g32485,g33459,I30995,I31466,g33318,g7909,g30038,g23253,I12103,
    I14668,I18734,g9681,g10040,g32555,g13028,g14536,g19860,g33458,g7519,g24361,
    g25557,g32570,g32712,g25210,g32914,g9914,g17613,g33918,g23236,g20500,
    g10621,g7567,g34677,g29365,g14252,g21175,g13664,g11252,I20318,g23952,
    g23351,g32907,I30641,g24049,I14896,g9820,g29960,g28885,g22881,g23821,
    g10564,g9462,I17401,g16075,g13597,g9413,g19659,g24048,g11576,I33064,I17989,
    g20004,g13484,g32567,g32594,g19658,g23264,g25286,g16623,g14127,g10183,
    g7586,g23516,g25039,g14183,I16770,g11609,g7660,g12903,g20613,g19422,g31817,
    g13312,g32941,g11608,g7659,g19644,g10509,g32519,I22031,g21387,g32675,g8388,
    g20273,g20106,g12563,g20605,g21422,I26409,I28458,g8216,g10851,I14069,
    g10872,g9601,g23422,g32518,I16328,g24106,g24605,I27391,g32637,g16920,
    I18265,g28153,g32935,g24463,I21769,g19402,g28314,g20033,g31823,g34329,
    g32883,g19411,g19527,g17710,g14764,g24033,g12845,g27990,g16853,g23542,
    g23021,I22576,g10213,g12899,g16589,g14082,g25169,g29955,g28950,g9060,
    g23913,I17392,g9460,g24795,g23342,g29970,I28199,g12898,g10405,I21959,
    g16588,g13929,I24334,g23614,g25410,g18829,I15732,g8741,g10047,I32812,
    g34588,g19503,g29878,g28421,g21607,g22999,g23607,g14205,g26654,g20514,
    g25222,g32501,g32729,g18828,g31631,I29221,g10311,I22419,g23905,g9739,
    g32577,I14730,g18946,g29171,g21274,g23274,g20507,g23530,g22998,g27832,
    g32728,g21346,g25015,g23662,g6977,g19714,I13240,g7275,g29967,g28946,g29994,
    g34531,g23565,g32438,g8883,g12440,g27573,g26667,g25556,I33176,g34887,g7174,
    g19979,I17970,g7374,g12861,g17651,g14868,g17672,g14720,g34676,g8217,I17471,
    g9390,g11214,g32906,g16285,g8466,g15732,g22449,g19597,g34654,I32766,g20541,
    g16305,g13346,g10350,g9501,g16809,g14387,g21409,g22897,g7239,g23409,g32622,
    g8365,g26851,g24789,g23309,g32566,g19741,g29079,g7380,g21408,g10152,g7591,
    g23408,g8055,g10396,g20325,g24359,g19067,g20920,g20535,g20434,g9704,g31816,
    g8133,I24089,g24535,g24358,g17505,g14899,g8774,g32653,I20216,g17717,g14937,
    g14386,g34222,I17166,g32138,g31233,g24121,I18888,g8396,g9250,g34587,I32671,
    g12997,g32636,I23998,g34577,g32415,g14405,g12170,g19695,g8538,g29977,
    g28920,I18066,g32852,g11235,g24641,g8509,g19526,g16630,g14142,I17901,
    g26814,g34543,g34359,g32963,g22148,I12000,g12871,g10378,g29353,g23537,
    g9568,g31842,g32664,g30569,I16345,g8418,g34569,g22646,g25465,g8290,g18903,
    g30568,g23283,g11991,g9485,g13414,g23492,g23303,g32576,g24134,g8093,g32484,
    g24029,g33424,g10113,g17811,g12925,g20506,I25750,g26823,g20028,g15371,
    g32554,g24506,g16194,g7750,g24028,I24784,g24265,g16712,g26841,g32609,
    g21381,g28779,g31830,g23982,I25369,g12181,g8181,I27253,g32608,g8381,g19689,
    g25117,g25000,g8685,g7440,g8700,g32921,g33713,g8397,g19688,g9626,g8021,
    g12735,g18990,g32745,g22896,g21012,g23840,g32799,g18898,g15566,g23390,
    g32813,I21810,g6820,g33705,g7666,g20649,g34391,g32798,I22353,g28380,g20240,
    I23387,g32973,g32424,g22716,g19795,g16675,g20648,g10881,g20903,g32805,
    g13082,g32674,g24648,g23148,g7528,g12859,g13107,I32659,g7648,g26615,g25432,
    g12950,g12708,g20604,g9683,g23522,g18832,g24604,g30578,g33460,I30998,
    g33686,g19885,g26720,g7655,I14602,g20770,I26508,g9778,g20563,g27996,g32732,
    g24770,g8631,g25230,g23314,g32934,g24981,g11849,g17582,g14768,g12996,
    g10027,g23483,g14198,g8301,g19763,g29976,g12844,g7410,g11398,g23862,g32692,
    g32761,I32648,g34371,g11652,g7674,g9661,g13141,g11374,g20767,g26340,g24953,
    g21326,g10710,I12300,g23948,g10204,g14204,g12155,g20633,g23904,g31837,
    g21252,g29669,g34275,g34047,g19480,g17603,g14993,g20191,g17742,g14971,
    g32539,g10081,I18168,g8441,g22857,g7235,g7343,g25007,g32538,g24718,g34580,
    g14786,g12471,g29195,g9484,g30983,g29657,g9439,g17681,g14735,g6840,g8673,
    g34983,I19756,g33455,g21183,g7693,g11833,g7134,g21397,g23847,g18061,g14800,
    I17609,g19431,I32089,g25116,g7548,I14158,g8669,g10090,g20573,I13699,g20247,
    g29893,g28755,g16622,g14104,g23509,g10182,g28620,g27679,g20389,g8058,
    g29382,g8531,g24389,g8458,g24045,g12902,g20612,g23508,I20870,g32771,g8743,
    g20388,g17297,g20324,g8890,g29713,g24099,g24388,g20701,g20777,g20534,
    g22317,g31623,g32683,g19670,g24534,g8505,g20272,g17239,I32071,g24098,
    g12738,g9616,g17504,g15021,g8011,g25340,g25035,g8734,g19734,g13106,g10897,
    g6954,g19930,g6810,g9527,g11812,I12314,g13463,g31822,g32515,g32882,g19694,
    g7908,g24032,g22626,g25517,g11033,g8500,g11371,g18911,g23452,g10026,g9546,
    g13033,g21205,g10212,g29939,g28857,I18180,g7518,I18117,g23912,g9970,g24061,
    g29093,g20766,g27980,g8080,g31853,g19502,g15674,g8480,I19796,g25193,g8713,
    g21051,g19618,g19443,g12895,g16585,g14075,g13514,g25523,g31836,g32441,
    g32584,g24360,g20447,g14149,g16609,g19469,I28336,g10620,g17737,g14810,
    g22856,g22995,g32759,g16200,g23350,g25006,g32725,I23330,g34522,g7933,
    g16608,g14116,g19468,g23820,g34952,g34351,g34174,g32758,g7521,g7050,g20629,
    g23152,g9516,g20451,g21396,g31616,I29214,g7231,g30063,g29015,g9771,I25552,
    g20911,g10369,g32744,g19677,g12490,g17512,g21413,g15585,g9299,I15788,
    g23413,g32849,g9547,g10368,g32940,g7379,g8400,g11724,g31809,g11325,g7543,
    g20071,g32848,g9892,g24071,g12889,I11632,g20591,g25781,g24510,g20776,
    g31808,g32652,g32804,g7289,g12888,g26614,g25426,g10133,g20147,g7835,g24147,
    g10229,g9478,g26607,g25382,g17499,g14885,g22989,g23929,I18293,g11344,g9015,
    g33838,g8806,g19410,g24825,g23204,g17498,g14688,g22988,g8183,g23020,g23928,
    g8608,g30021,g28994,g33665,g19479,g19666,g17188,g6782,g25264,g16692,g14170,
    g25790,g29705,g25137,I13094,g17056,g30300,g11291,I32591,g34287,g23046,
    g32962,I14823,g19478,g24996,g17611,g14822,g9907,g13173,g12377,g30293,
    I16698,I31724,g9959,g8977,g24367,g24394,g32500,g9517,g9690,g23787,g29170,
    g32833,g18957,g21282,g16214,I32950,g23282,g7541,g10627,I13968,g34320,
    g34119,g27089,g23302,g25209,g19580,g30593,I31500,g6998,g22199,g34530,
    g10112,g7132,g12546,g10050,g27088,g26694,g34346,g34162,g25208,g7153,g7680,
    g8451,g22198,g22529,g19549,I32059,g15799,g13110,g13506,g10808,g12088,g7701,
    g20446,g9915,g12860,g22528,g23769,g22330,g25542,g7802,g20059,g32613,g8146,
    g10096,g20025,g8346,g24059,g33454,g24025,g9214,g17529,g15039,g20540,g16646,
    g12497,g30292,g28736,g10615,g23768,g20058,g24540,g33712,g32947,g19531,
    g24058,g22869,g17528,g14940,g7558,I12041,g32605,g8696,g19264,g22868,g11927,
    g10207,g23881,g10857,g32812,g32463,g19676,g19685,g31239,g29916,g25274,
    g24044,g16771,g14018,g19373,g26575,g25268,g10428,g32951,g32972,g16235,
    g32033,g30929,g8508,g19654,g9402,g9824,g8944,g8240,g18661,g18895,g19800,
    g21662,g24377,g24120,g23027,g32795,g25034,g23695,g23299,g17709,g14761,
    g33382,g8443,g20146,g20738,g20562,g9590,g21249,g11290,g24146,g23249,g20699,
    g16515,g13486,g10504,g11981,g9657,g12968,g17471,g25153,g8316,g17087,g23482,
    g32514,g24699,g23047,g21248,g14504,g12361,g19762,g23248,g19964,g20698,
    g27527,g25409,g34575,g32507,g9556,g8565,g21204,g33637,g29177,g34711,g12870,
    g25136,g34327,g34108,g10129,g9064,g8681,g10002,g10057,g9899,g34367,g7262,
    g24366,g20632,g8697,g24374,g19543,g30303,g28786,g8914,g17602,g14962,g12867,
    g10375,g12894,g16584,g13920,g17774,g14902,g23647,g18889,g18980,g32541,
    g10323,g23945,g16206,g24481,g23356,g32473,I31463,g26840,g20661,g21380,
    g10533,g20547,g23999,g32789,g18888,g23380,g20619,g33729,g19569,g16725,
    g13963,g13521,g11357,g22994,g32788,g32724,g19747,g23233,g21182,g6789,
    g11832,g23182,g21389,g20715,g32829,g32920,g32535,g25327,g22161,g32434,
    I21258,g25109,g12818,g20551,g20572,g15833,g9194,g32828,g18931,g32946,
    g10232,I17276,g7285,g11861,g22919,g14232,g11083,g9731,g23331,g20905,g34397,
    g19751,g16044,g24298,g9489,g19772,g25283,I22177,g23449,g26483,g9557,g24127,
    g13045,g10261,g23897,g11324,g23448,g23961,g32682,g24490,g34192,g33921,
    g16652,g13892,g23505,g26326,g24872,g20385,g19416,g20103,g7424,g24376,
    g24385,g7809,g24103,g23026,g24980,I12117,g24095,g26702,g17599,g14794,
    g25174,g23890,g28696,g31653,g6991,I14939,g20671,g14844,g27018,g31138,
    g29778,g32760,g17086,g7523,g19579,g22159,g29941,g28900,g13140,g7643,g12018,
    g9538,g34553,g10499,g32506,I21288,g29092,g34949,g34326,g34091,g13061,
    I18479,g31852,g6959,g30040,g29025,g19586,I12123,g27402,g34536,g30307,
    g23433,g34475,g24426,g8479,g20190,g22144,I24038,g10080,g34388,g8840,g9212,
    g12866,g21343,g8390,g32927,g14432,g12311,g17680,g14889,g17144,g14085,
    g26634,g25317,g7926,g20546,g20089,g23971,I26378,g19720,g20211,g24089,
    g27597,g26745,g21369,g12077,g32649,g25553,g20088,g9229,g14753,g24088,
    g19493,g24024,g14342,g12163,g34673,g31609,g10031,g32648,g32491,g32903,
    g25326,g10199,g16605,g13955,g11472,g7918,g31608,g29653,g20497,g32604,
    g34062,g33711,g32755,I30959,g11911,g10022,g16812,g21412,g32770,g12180,
    g32563,g13246,g20700,g20659,g20625,g24126,g24625,g23135,g24987,g8954,
    g31799,g23896,g25564,g22312,g8363,g18894,g31813,g21228,g33799,g33299,
    g10365,g22224,g33813,g19517,g23228,g29906,g28793,g29348,g28194,g10960,
    g23011,g31798,g32767,g32794,g11147,g8417,g11754,g25183,g32899,g7534,g31805,
    g16514,g14139,g12885,g22495,g17308,g14876,g23582,I22729,g32633,g32898,
    g9620,g19362,g16072,g7927,g34574,g32719,g18979,g19523,g24060,g33934,g10708,
    g7836,g20197,g21379,g34311,g34097,g22985,g32718,g32521,I13597,g23925,
    g18978,g21050,g20527,g11367,g32832,g23378,g33761,g24527,g7903,g17687,
    g15042,I31604,g10043,g7513,g26731,g25470,g29333,g28167,g16473,g13977,
    g32861,g9842,g23944,g32573,g31013,g29679,g25213,g23293,g19437,g20503,g9298,
    g28598,g27717,g32926,g7178,g7436,g29963,g28931,g16724,g14079,g22842,g19875,
    g23681,g32612,g16325,g18877,g25452,g25047,g32099,g31009,g18216,g34820,
    g20714,g20450,g23429,g32701,g7335,g7831,g32777,g32534,g12721,g20707,g21428,
    g20910,g23793,g12054,g7690,g17392,g14924,g19600,g10337,g24819,g19781,
    g17489,g20496,g7805,g25051,g25072,g32462,g24979,g21690,g22830,g19952,
    g24055,g7749,g19351,g23549,g20070,g16173,g20978,g24111,g28656,g9708,g24070,
    g24978,g34691,g29312,g28877,g20590,g22544,g19589,g22865,g23548,g8778,
    g29115,g7947,g24986,g9252,g23504,g13902,g11389,g13301,g18917,g19790,g20384,
    g9958,g29921,g28864,g13120,g24384,g25820,g20067,g32766,g6955,g29745,g28500,
    g24067,g24094,g11562,g17713,g12947,g8075,g32871,g30020,g22189,g9829,g12839,
    g6814,g12930,g12347,g7873,g26743,g25476,g26827,g34583,g21057,g10079,g24150,
    g23057,g9911,g7495,g14545,g12768,g7437,g17610,g15008,g12838,g10353,g23128,
    g16486,g10078,g24019,g17189,g14708,g23245,g26769,g8526,g19208,g21299,
    g30113,g29154,g9733,g10086,g23323,g9974,g17124,g14051,g26803,g12487,g20526,
    g24526,g19542,g30302,g28924,g7752,g18102,g8439,g9073,g32629,g27277,g30105,
    g7917,g27279,g26330,g32472,g10159,g34827,g10532,g32628,g32911,g15344,
    g14851,g10158,g11403,g11547,g20917,g19905,g18876,g18885,g25046,g23729,
    g6993,g10295,g13715,g27038,g25932,g32591,g23995,g32776,g32785,g19565,
    g24077,g20706,g23880,g20597,g32754,g7932,g25282,g27187,g7296,g23512,g8616,
    g20923,g27975,g32859,g32825,g32950,g26710,g18660,g20624,g22455,g12975,
    g12752,g7532,g11171,g32858,g33744,g7553,g8404,g31849,g8647,g14631,g12239,
    g19409,g20102,g20157,g12937,g12419,g28669,g27705,g24619,g8764,g22201,
    g24102,g23445,g31848,g18916,g24157,g32844,g9898,g33848,g33261,g28260,
    g27703,g17617,g7885,g18550,g25768,g25803,g24798,g31141,g12224,I26960,
    g22075,g18314,g33652,g33393,g18287,g27410,g16633,g30248,g28743,g34482,
    g34405,g23498,g20234,g28489,g27010,g26356,g15581,g18307,g29771,g28322,
    g30003,g28149,g34710,g16191,g22623,g19337,g21989,g30204,g28670,g13671,
    g26826,g24907,g27666,g26865,I31246,g18721,g15138,g22037,g25881,g26380,
    g19572,g33263,g18596,g32420,g31127,g28488,g27969,g27363,g23056,g16052,
    g27217,g26236,g29683,g18243,g33332,g32217,I17692,g14988,g21988,g26090,
    g21924,g28558,g18431,g26233,I31071,g26182,g26651,g22707,g12015,g34081,
    g33706,g27486,g31962,g24763,g17569,g33406,g32355,g18269,g15069,g33361,
    g32257,g15903,g13796,g18773,I31147,g18341,g29515,g28888,g29882,g18268,
    g29991,g29179,g21753,g31500,g29802,g18156,g18655,g15106,g33500,I31196,
    I31197,g24660,g22648,g33833,g33093,g32203,g18180,g26513,g19501,g17418,
    g14407,I27409,g34999,g18670,g34380,g34158,g25482,I24597,g32044,g31483,
    I24684,g16612,g21736,g11546,g21887,g15101,g30233,g28720,g18734,I31151,
    g16324,g13657,I31172,g18335,g16701,g22589,g19267,g32281,g31257,g34182,
    g28255,g16534,g28679,g27572,g11024,g16098,I13937,g18993,g11224,g24550,
    g32301,g31276,g14643,g11998,g12023,g24314,g22588,g21843,g32120,g24287,
    g28124,g27368,g15794,g18667,g18694,g12179,g24307,g29584,g27178,g21764,
    g11497,g18131,g29206,I27528,I27529,g13497,g28686,g27574,g32146,g17321,
    g27421,g24721,g17488,g22119,g21869,g27186,g26195,g31273,g30143,g34513,
    g21960,g27676,g26377,g27685,g13032,g15633,g33106,g32408,g18487,g27373,
    g29759,g28308,g22118,g32290,g31267,g11126,g12186,g28267,g17401,g13143,
    g21868,g18619,g18502,g22022,g34961,g12953,g18557,g18210,g29758,g28306,
    g17119,g33463,I31011,I31012,I31227,g18618,g18443,g24773,g22832,g21709,
    g18279,g30026,g28476,g33371,g32280,g30212,g28687,g16766,g26387,g24813,
    g27334,g12539,g34212,g28219,g21708,g15049,g18278,I16111,g11409,g11381,
    g26148,g25357,g16871,g29345,g22053,g23471,g20148,g26097,g18469,g24670,
    g33795,g33138,g28218,g27768,g29940,g26104,g18286,g22900,g17137,g26218,
    g15861,g8690,g27964,g25956,g18468,g25331,I24508,g18306,g15074,g12762,
    g22036,g25449,g13060,g31514,g32403,g31117,g27216,g33514,I31266,I31267,
    g22101,g24930,g29652,g29804,g17809,I31281,g28160,g26309,g15612,g22680,
    g18815,g30149,g28605,g25961,g25199,I27381,g33507,I31231,I31232,I31301,
    g20131,g15170,g15701,g10705,g18601,g13411,g11834,g18187,g18677,g14610,
    g28455,g27289,g33421,g32374,g21810,g17177,g21774,g29332,g29107,g23657,
    g19401,g28617,g27533,g21955,g23774,g14867,g22064,g15162,I24600,I31146,
    g22929,g34104,g27117,g21879,g34811,g14165,g21970,g18143,g24502,g23428,
    g28201,g27499,g19536,g19948,g17515,g29962,g23616,g21878,I16695,g12523,
    g12463,g32127,g31541,g22536,g24618,g22625,g26229,g33473,I31061,I31062,
    g18169,g21886,g27568,g18791,g31789,g30201,g28467,g26993,g28494,g27973,
    g33789,g33159,g21792,g16591,g22009,g22665,g17174,g18168,g18410,g21967,
    g21994,g31788,g33724,g14145,g32376,g19564,g17175,g33359,g32252,g25149,
    g14030,g17693,g22008,g32103,g24286,g18479,g18666,g33829,g33240,g18363,
    g32095,g18217,g15063,g33434,g32239,g24306,g33358,g32249,g25148,g16867,
    g11496,g15871,g18478,g30133,g28591,g33828,g33090,g28352,g11111,g14875,
    g34133,g21919,g15144,g30229,g28716,g25104,g16800,g11978,g26310,g23919,
    g32181,g31020,g33121,g18486,g27230,g25906,g27293,g9972,g29613,g28208,
    g28266,g23748,g19062,g33344,g32228,g14218,g21918,g30228,g28715,g26379,
    g19904,g18556,g25971,g24187,g34228,g30011,g29183,g27265,g26785,I31226,
    g16844,g18580,g26050,g27416,g26314,g26378,g19576,g13384,g11804,g29605,
    g18223,g27992,g26800,g22074,g27391,g24143,g25368,g27510,g7764,g32190,
    g26096,g29951,g18110,g34310,g14003,g25850,g15911,g28588,g27489,g28524,
    I31127,g18321,g24884,I24051,g30925,g29908,g21817,g11019,g18179,g13019,
    g18531,g30112,g28566,g28477,g27966,g33760,g33143,g24410,g32089,g27261,
    g25229,g30050,g22545,g29795,g28344,g18178,g18740,g26857,g25062,g25049,
    g34050,g21977,g22092,g23532,g19400,g23901,g13095,g16025,g33506,I24530,
    g32088,g27241,g24666,g22518,g12982,g21783,I31297,g24217,g18186,g15785,
    g18676,g18685,g10800,g18373,g29514,g24015,g19540,g30096,g28546,g22637,
    g19363,g17176,g34742,g28616,g27532,g18654,g16203,g28313,g27231,g27116,
    I27509,g21823,g27615,g26789,g18800,g15859,I31181,g18417,g24556,g28285,
    g34681,I27508,g15858,g27041,g32126,g18334,g27275,g25945,g19756,g33927,
    g33094,g28254,g27395,g27430,g34857,g10822,g24223,g27493,g16957,g25959,
    g30730,g26346,g25925,g24990,g28466,g27960,g25112,g21966,g18762,g25050,
    g13056,g20084,g11591,g32339,g31474,g31240,g14793,g15968,g34765,g27340,
    g27035,g26348,g18423,g12851,g29789,g28270,g32338,g31466,g33491,I31152,
    g33903,g33447,g24922,g26129,g24321,g16699,g27684,g26386,g28642,g27555,
    g18587,g25096,g23778,g29788,g28335,g26128,g14589,g10586,g10569,g29535,
    I31211,g27517,g18909,g16226,g32197,g31144,g18543,g26323,g24186,g14588,
    g11957,g11974,g24676,I16721,g12589,g12525,g18117,g16427,g25802,g22083,
    g32411,g31119,g23023,g19691,g24654,g28630,g27544,g29344,g29168,g18569,
    g30002,g28481,g27130,g30057,g29144,g22622,g19336,g18568,g18747,g25765,
    g24989,g24973,g27362,g26080,g31990,g31772,g33899,g18242,g10616,g27523,
    g30245,g28733,I31126,g26232,g33898,g33419,g21816,g18123,g18814,g33719,
    g33141,g24762,g10704,g34533,g34318,g18751,g18807,g21976,g21985,g15902,
    g18772,g28555,g27429,g33718,g33147,g8679,g28454,g26976,g33521,I31302,
    g18974,g26261,g24688,g32315,g31306,g24423,g21752,I31296,g18639,g28570,
    g27456,g28712,g27590,g21954,g27222,g29760,g28309,g33832,g33088,g18230,
    g14506,g27494,g17139,g18293,I18620,g15738,g18638,g27437,g33440,g32250,
    g32055,g10999,g17138,g18265,g25129,g17682,g15699,g30232,g28719,g32111,
    g18416,g25057,g23275,g32070,g10967,g33861,g33271,g28239,g27135,g25128,
    g17636,g10829,g11916,g33247,g32130,g28567,g27347,g18992,g18391,g24908,
    I24075,g28238,g27133,g21842,g18510,g30261,g28772,g23392,g24569,g25323,
    g31324,g30171,g33099,g32395,g13287,g27600,g26755,g10733,g18579,g31777,
    g33701,g33162,g24747,g17510,g32067,g21559,g16236,g31272,g30117,I16618,
    g12341,g12293,g15632,g28185,g27026,g18578,g25775,g23424,g27351,g27372,
    g19768,g14874,g16671,g21558,g15904,g27821,g32150,g28154,g18586,g29649,
    g33462,I31006,I31007,g21830,g26611,g24935,g16260,g10665,g28637,g22399,
    g18442,g32019,g30579,g24772,g16287,g29648,g27264,g25941,g22115,g27137,
    g21865,g31140,g32196,g27587,g13942,g24639,g32018,g26271,g29604,g30316,
    g29199,g21713,g31288,g24230,g13156,g18116,g24293,g18615,g22052,I13862,
    g24638,g29770,g28320,g16190,g14626,g29563,I31202,g13888,g18720,g15137,
    g26753,g16024,I31257,g25880,g14555,g12521,g12356,g12307,I16671,g24416,
    g16520,g21705,g30056,g29165,g18275,g15070,g26145,g11962,I31111,g18430,
    g18746,g27209,g26213,g32402,g18493,g33871,g33281,g30080,g28215,g26650,
    g10796,g16211,g27208,g18465,g29767,g28317,g29794,g28342,g21188,g33360,
    g32253,g18237,g29845,g28375,g23188,g13994,I16143,g11491,g11445,g28439,
    g27273,g18340,g29899,g28428,g29990,g29007,g21939,g25831,g15784,g18806,
    g18684,g26393,g19467,g14567,g10568,g10552,g24835,g8720,g29633,I31067,
    g24014,g15103,g34753,g21938,g18142,g34342,g34103,g30145,g28603,g30031,
    g29071,g27614,g32256,g31249,g18517,g27436,g30199,g28664,g29718,g28512,
    g29521,g16700,g31220,g30273,g33472,I31056,I31057,g16126,g28284,g10675,
    g25989,g25258,g27073,g26281,g30198,g28662,g32300,g31274,g14185,g25056,
    g28304,g27226,g33911,g33137,g34198,g26161,g34529,g34306,g21875,g25988,
    g25924,g24976,g27346,g34528,g34305,g17692,g18130,g34696,g18193,g22013,
    g32157,g34393,g34189,g26259,g24430,g18362,g23218,g20200,g29861,g28390,
    g29573,g33071,g21837,g34764,g22329,g11940,g10883,g18165,g23837,g18523,
    g26087,g27034,g26328,g13306,g31776,g34365,g34149,g26258,g19651,g16119,
    g33785,g33100,g29926,g34869,g28139,g27337,g22005,g31147,g12286,g28653,
    g13038,g27292,g29612,g27875,g24465,g22538,g14035,g27153,g33355,g32243,
    g29324,g29078,g34868,g7396,g25031,g20675,g30161,g28614,g18475,g12853,
    g33859,g26244,g29534,g28965,g33370,g32279,g24983,g23217,g27409,g16855,
    g28415,g27250,g24684,g28333,g27239,g33858,g33268,g34709,g18222,g10501,
    g16870,g27136,g27408,g27635,g21915,g30225,g28705,g31151,g18437,g24142,
    I31001,g31996,g31779,g34225,I31077,g26602,g30258,g28751,g11937,g15860,
    g23201,g14027,g33844,g33257,g33367,g32271,I31256,g18703,g22100,g18347,
    g19717,g14438,g10726,g30043,g29106,g18253,g25132,g30244,g28732,g26171,
    g15700,g18600,g20193,g15578,g18781,g28585,g27063,g24193,g28484,g10290,
    I26972,g33420,g32373,g30069,g29175,g29766,g28316,g18236,g15065,g21782,
    g17771,g13288,g20165,g34069,g21984,I31102,g26994,g26226,g27474,g28554,
    g27426,I31157,g18351,g18372,g24523,g22318,g32314,g31304,g29871,g28400,
    g33446,g32385,g26166,g16707,g21419,g16681,g32287,g34774,g34695,g18175,
    g18821,g15168,g34931,g27327,g13077,g16202,g28312,g27828,g28200,g27652,
    g32307,g31291,g14566,g10566,g10551,g32085,g27253,I31066,g29360,g27364,
    g21822,g22515,g12981,g22991,g27537,g28115,g27354,g31540,g29904,g25087,
    g17307,g32054,g10890,g24475,g7685,g18264,g18790,g18137,I27513,g18516,
    g34337,g34095,g24727,g13300,g34171,g33925,g16590,g24222,g16986,g27303,
    g11996,g11223,g25043,g20733,g32269,g31253,g21853,g28799,g27445,g26079,
    g34967,g28813,g29629,g28211,g32341,g31472,g31281,g30106,g15870,g26078,
    g32156,g25069,g23296,g24703,g17592,g31301,g30170,g18209,g29628,g27924,
    g33902,g33085,g21836,g31120,g32180,g23836,g26086,g28674,g27569,g13321,
    g25068,g17574,g25955,g24720,g30919,g29898,g18208,g16801,g16735,g23401,
    g25879,g11135,g24600,g22591,g25970,g31146,g12285,g30010,g29035,g30918,
    g32335,g11178,g11740,g8769,g18542,I18803,g18453,g29591,g28552,g29785,
    g28332,g31290,g29734,g22114,g26159,g26125,g21864,g34079,g33703,g22082,
    g27390,g26977,g30599,g22107,g30078,g28526,g21749,g26158,I18716,g26783,
    g25037,I31287,g18614,g28692,g27578,g28761,g34078,g33699,g18436,g25967,
    g30598,g14585,g29859,g28388,I31307,I31076,g30086,g28536,g21748,g15089,
    g15707,g15819,g18607,g18320,g24790,g21276,g17625,g21285,g7857,g26295,
    g29858,g28387,g21704,g22849,g33366,g32268,g27522,g24401,g15818,g18530,
    g25459,I24582,g18593,g18346,g19716,g12100,g21809,g23254,g20056,g28214,
    g27731,g15111,g22848,g19449,g18122,g15052,g23900,g34322,g14188,g14608,
    g12638,g12476,g12429,g15978,g18565,g26336,g10307,g30125,g28581,g18464,
    g21808,g29844,g28374,g34532,g34314,g15590,g29367,g28539,g10921,g27483,
    g30158,g28613,g33403,g32352,g24422,I31341,g32278,g27553,g26293,g18641,
    g18797,g25079,g21011,I31156,g18292,g16706,g31226,g30282,g32286,g34561,
    g34368,g16597,g18153,g27326,g12048,g25078,g23298,g31481,g29768,g32039,
    g31476,g33715,g33135,g32306,g31289,g34295,g34057,g33481,I31101,g22135,
    g27536,g18409,g27040,g25086,g13941,g21733,g10674,g18136,g18408,g18635,
    g24726,g15965,g27252,g26733,g24913,g21874,g25817,g24807,g32187,g30672,
    g26289,g24436,g25159,g10732,g22049,g25125,g20187,g27564,g26305,g25901,
    g24853,g26023,g9528,I31131,g34966,g31490,g29786,g10934,g24607,g25977,
    g25236,g26288,g33490,g19681,g24320,g28235,g26571,g10472,g23166,g13959,
    g20196,g22048,g26308,g29203,I27514,g18164,g28683,g27876,g32143,g31784,
    g30176,g34364,g34048,g33784,g33107,g24952,g31297,g30144,g27183,g33376,
    g32294,g27673,g25769,g22004,g23008,g33889,g33303,g11123,g24464,I24027,
    g16885,g32169,g31014,g18575,g18474,g29902,g28430,g30289,g28884,g29377,
    g28132,g13807,g18711,g15136,g32168,g30597,g32410,g27469,g13974,g18327,
    g24797,g22872,g30023,g21712,I24482,g18109,g27508,g16763,g27634,g26805,
    g34309,g13947,g21914,g24292,g30224,g28704,g18537,I24710,g34224,g30308,
    g29178,g22106,I24552,g29645,I24003,I18568,g27225,g18108,g14207,g21907,
    I31286,g15077,g24409,g25966,I31306,g13265,g18283,g13296,g18606,g18492,
    g18303,g24408,g23989,g24635,g19874,g34495,g34274,g22033,g27213,g18750,
    g15145,g31520,g29879,I31187,g33520,g18982,g18381,g34687,g14181,g21941,
    g26842,I27429,g27452,g21382,g29632,g28899,g31211,g34752,g18174,g27311,
    g12431,g18796,g28725,g27596,g32084,g10948,g32110,g16596,g25571,I24694,
    I24695,g33860,g33270,g32321,g27613,g16243,g29661,g29547,g29895,g28107,
    g27970,g10683,g32179,g31748,g21935,g18390,g31497,g33497,I31182,g20109,
    g17954,g24327,g21883,g32178,g31747,g15876,g13512,g11116,g20108,g15508,
    g34842,g34762,g18192,g22012,g26544,I27504,g25816,g33700,g33148,g33126,
    g31987,g31767,g29551,g29572,g26713,g25447,I31217,g34489,g34421,g24283,
    g18522,g27350,g18663,g24606,g25976,g24303,g16670,g27820,g34525,g34297,
    g28141,g11797,g34488,g34417,g27282,g13493,g25374,I24527,g31943,I24505,
    g21729,g26610,g33339,g32221,g33943,g33384,g31296,g30119,g34558,g34353,
    g16734,g23577,g19444,g18483,g24750,g17662,g32334,g31375,g21728,g33338,
    g32220,g28263,g23747,g16930,g23439,g13771,g11035,g18553,g13035,g26270,
    g31969,g29784,g28331,g26124,g22920,g19764,g16667,g20174,g29376,g14002,
    g27413,g34865,g16965,g18949,g31968,g31757,g18326,g24796,g11142,g27691,
    g25778,I18713,g29354,I27533,g18536,g23349,g13662,g22121,g29888,g28418,
    g33855,g33265,g14206,g21906,g18702,g15133,g21348,g18757,g31527,g23083,
    g16076,g23348,g15570,g15076,g33870,g33280,g33411,g32361,g33527,I31331,
    I31332,g26294,I31321,g16619,g30042,g29142,g18252,g18621,g25559,g13004,
    g30255,g28748,g25488,I24603,g28833,g16618,g34679,g14093,g18564,g30188,
    g28644,g24192,g30124,g28580,g16279,g34678,g31503,I31186,g33503,I31212,
    g24663,g16621,g33867,g33277,g14637,g34686,g34494,g13523,g18183,g18673,
    g25865,g25545,g18397,g30030,g29198,g30267,g28776,g33450,g32266,g22760,
    g22134,g27113,g32242,g31245,g18509,g22029,g31707,g30081,g34065,g33707,
    g33174,g18933,g16237,g33910,g33134,g24553,g22983,g26160,g28273,g27927,
    g7696,g18508,g22028,g27302,g18634,g21333,g23415,g20077,g27357,g25042,
    g23262,g31496,g33818,g33236,g24949,g23796,g33496,I31176,I31177,g19461,
    g11708,g27105,g24326,g30219,g28698,g17134,g21852,g15839,g34875,g28812,
    g26972,g33111,g34219,g25985,g19145,g24536,g19516,g29860,g28389,g17506,
    g14505,g25124,g15694,g15838,g21963,g24702,g17464,g34218,g24757,g31986,
    g31766,g19736,g12136,g24904,g11761,g28234,g27877,g32293,I31216,g25939,
    g24583,g26277,g18213,g32265,g25030,g23251,g25938,g25093,g31067,g29484,
    g24564,g23198,g29625,g28514,g29197,g19393,g16884,g18574,g23484,g20160,
    g18452,g18205,g31150,g23554,g20390,I31117,g18311,g33801,g33437,g24673,
    g22659,g33735,g33118,g33877,g33287,g30915,g29886,g29943,g7834,g16666,
    g25875,g31019,g29481,I18765,g29644,g28216,g29338,g29145,g30277,g28817,
    g13063,g31018,g29480,g32014,g29969,g30075,g28525,g26155,g14221,g21921,
    g26822,g24841,I31242,g18592,g23921,g18756,g34075,g33692,g31526,g22521,
    g24634,g22634,g30595,g33526,I31326,I31327,g29968,g21745,g18780,g12027,
    g14613,g10602,g10585,g27249,g25929,g21799,g29855,g17770,g21813,g23799,
    g14911,g27482,g15815,g28541,g27403,g10947,g18350,g33402,g32351,g29870,
    g29527,g28945,g27710,g26422,g21798,g34782,g18820,g15166,g26853,g28789,
    g27440,g21973,g32116,g27204,g33866,g33276,g22899,g19486,g21805,g22990,
    g19555,g18152,g25915,g24926,g32041,g13913,g18396,g22633,g19359,g18731,
    g15140,g30266,g28775,g28535,g15937,g11950,g25201,g12346,g22191,g16179,
    g29867,g29894,g19069,g21732,g16531,g13542,g21934,g18413,g24912,g23687,
    g26119,g11944,g24311,g16178,g18691,g15884,g33689,g33144,g32340,g31468,
    g29581,g28462,g32035,g31280,g29717,g17191,g17719,g14675,g21761,g29315,
    g29188,g27999,g26200,g26864,g26022,g25271,g13436,g18405,g31300,g30148,
    g30167,g28622,g30194,g28651,g30589,I24690,I24549,g26749,g24494,g27090,
    g29202,g25782,g32142,g13320,g26313,g12645,g28291,g29979,g23655,g26082,
    g22861,g19792,g27651,g22448,g34524,g33102,g32399,g26276,g26285,g34401,
    g34199,g26344,g22045,g18583,g29590,g26254,g31066,g29483,g31231,g30290,
    g29986,g28468,g22099,g27932,g25944,g27331,g30118,g28574,g24820,g13944,
    g26808,g25521,g16762,g20152,g11545,g22534,g28179,g22098,g32193,g30732,
    I31116,g24846,I24018,g26101,g33876,g33286,g33885,g33296,g26177,g18113,
    g18787,g15158,g32165,g31669,g24731,I31041,g18282,g34748,g27505,g27404,
    g31763,g30127,g18302,g33511,I31251,I31252,g18357,g19545,g29877,g28405,
    g15110,g18105,g10724,g22032,g30254,g28747,g18743,g27212,I31237,g21771,
    g10828,g18640,g18769,g15151,g22061,g30101,g28551,g30177,g28631,g29526,
    g28938,g17140,g26630,g34560,g34366,g18768,g18803,g15161,g31480,I31142,
    g33480,I31096,I31097,g24929,g23751,g22871,g27723,g26512,g15654,g31314,
    g30183,g28240,g27356,g27149,g30064,g28517,I18762,g27433,g27387,g15936,
    g25285,g22152,g29866,g27148,g21882,g21991,g26485,g24968,g23991,g19209,
    g27097,g25867,g33721,g33163,g19656,g27104,g16751,g13155,g16807,g27646,
    g13094,g25900,g24390,g34874,g23407,g9295,g33243,g32124,g28563,g25466,
    g23574,g19680,g12028,g33431,g16639,g26712,g24508,I17741,g18662,g15126,
    g32175,g31709,g30166,g28621,g30009,g29034,g24302,g15124,g16638,g33269,
    g31970,g34665,g21289,g18890,g13492,g27369,g25894,g24743,g22708,g30008,
    g29191,g18249,g33942,g33383,g33341,g32223,g18482,g10755,g29688,g29624,
    g28491,g14028,g18248,g15067,g16841,g18710,g15135,g34476,g34399,g34485,
    g34411,g18552,g24640,g24769,g19619,g19631,g16093,g18204,I31222,g27412,
    g34555,g34349,g18779,g22071,g24803,g22901,g33734,I31593,g30914,g29873,
    g21759,g15117,g23725,g14772,g18778,g25874,g11118,g27229,g31993,g31774,
    g21758,g26176,g26092,g18786,g15156,g27228,g24881,I24048,I31347,g22859,
    g26154,g30239,g28728,g17785,g13341,g25166,g31131,g18647,g34074,g33685,
    g30594,g18356,g29876,g28404,g29885,g28416,g21744,g30238,g28727,g34567,
    g34377,I31600,g28440,g27274,g18826,g18380,g19571,g33487,I31132,g22172,
    g29854,g21849,g21940,I31236,g15814,g31502,g28573,g25485,g33502,I31206,
    I31207,g29511,g31210,I31351,g18233,g28247,g27147,g21848,g15807,g18182,
    g27310,g26574,g18651,g15102,g18672,g15127,g34382,g34167,g30185,g28640,
    g34519,g34293,g17151,g21804,g34185,g27627,g13266,g25570,I24689,g27959,
    g25948,g28612,g27524,g30154,g28611,g28324,g24482,g31278,g29716,g34518,
    g34292,g32274,g31256,g27050,g25789,g27958,g25950,g25907,g24799,g24710,
    g22679,g27378,g26089,I31137,g18331,I27364,g24552,g22487,g33469,I31042,
    g28251,g27826,g30935,g28272,g27721,g31286,g30159,g32122,g18513,g21332,
    g18449,g12852,g27386,g19752,g33468,I31036,I31037,g15841,g25567,I24674,
    I24675,g27096,g18448,g29550,g28990,g32034,g14124,g25238,g12466,g16806,
    g29314,g29005,g22059,g21962,g18505,g21361,g7869,g22025,g18404,g24786,
    g33815,g33449,g32292,g31269,g10898,g18717,g22058,g31187,g32153,g24647,
    g19903,g33677,g31975,g31761,g13252,g11561,g11511,g11469,g18212,g29596,
    g27823,g24945,g23183,g10719,g16517,g21833,g15096,g30215,g28690,g32409,
    g14719,g34215,g30577,g26267,g24577,g25518,I24625,g27428,g13564,g22044,
    g26304,g31143,g29506,I24709,I31021,g24998,g17412,g12730,g27765,g24651,
    g24672,g19534,g14832,g29773,g28203,g27690,g25784,g16193,g27549,g31169,
    g11397,g18723,g25883,g13728,g28360,g27401,g22120,g33884,g33295,g15116,
    g18149,g27548,g31168,g32164,g30733,g18433,g33410,g32360,g18387,g24331,
    g30083,g28533,g13509,g27504,g18620,g18148,g21947,g30284,g28852,g34083,
    g33714,g34348,g34125,g33479,I31091,I31092,g34284,g34046,g21605,g13005,
    I31346,g33363,g32262,g13508,g18104,g18811,g18646,I31122,g14612,g11971,
    g11993,g31478,g29764,g8234,g31015,g29476,g18343,g12847,g24897,I24064,
    g29839,g30566,g26247,g33478,I31086,I31087,g24961,g23193,g21812,g17146,
    g34566,g34376,g28451,g27283,g16222,g31486,g29777,g32327,g31319,g29667,
    g29838,g27129,g33486,g32109,g21951,g26852,g24975,g24958,g21972,g15152,
    g27057,g19610,g16069,g18369,g12848,g24717,g22684,g27128,g28246,I31292,
    g32108,g30139,g28596,g18368,g34139,g16703,g22632,g19356,g31223,g21795,
    g32283,g31259,g27323,g26268,g30138,g28595,g27299,g26546,g29619,g32303,
    g27550,g34138,g11047,g18412,I31136,g11205,g13047,g27298,g26573,g29618,
    g28870,g19383,g16893,g34415,g34207,g18133,g15055,g23514,g20149,g26484,
    g24946,g33110,g13912,g9984,g24723,g17490,g31321,g30146,g18229,g33922,
    g33448,g14061,g33531,I31352,g18228,g24387,g26312,g34963,g32174,g31708,
    g16321,g16304,g28151,g18716,g31186,g33186,g32037,g24646,g22640,g33676,
    g33125,g33373,g32288,g16516,g27697,g25785,g18582,g27995,g26809,g31654,
    g29325,g30576,g22127,g24705,g34484,g34407,g18310,g29601,g31936,g33417,
    g32371,g21789,g26799,g25247,g29975,g28986,g34554,g34347,g18627,g15093,
    g15863,g13762,g18379,g30200,g28665,g21788,g33334,g32219,g18112,g16422,
    g13627,g23724,g14767,g18378,g22103,g15164,g21829,g29937,g13044,g14220,
    g21920,g23920,g22095,g16208,g25963,g28318,g27233,g18386,g30921,g29900,
    g28227,g21828,g15703,g17784,g18603,g21946,g18742,g33423,g32225,g29884,
    g34745,g27316,g24228,g18681,g24011,g32326,g31317,g29666,g28980,g17181,
    g16614,g17671,g29363,g23682,g16970,g18802,g18429,g32040,g14122,g24716,
    g15935,I24680,g33909,g33131,g34184,g18730,g15821,g27988,g26781,g18793,
    g18428,g24582,g33908,g33092,g28281,g16593,g12924,g27432,g13020,g18765,
    g28301,g27224,g24310,g16122,g18690,g15130,g28739,g18549,g11046,g25921,
    g24936,g13046,g26207,g24627,g29580,g28519,g21760,g20112,g13540,g31242,
    g29373,g22089,g27461,g33242,g32123,g18548,g15873,g28645,g27556,I31192,
    g27342,g12592,g24378,g16641,g27145,g14121,g22088,g18504,g22024,g31123,
    g32183,g19266,g33814,g33098,g28290,g23780,g32397,g31068,g13282,g27650,
    g29110,g12687,g25973,g18317,g12846,g33807,g33112,g31974,g31760,g29321,
    g29033,g33639,g33386,g26241,g34214,g29531,g31230,g30285,g18129,g30207,
    g28680,g16635,g27696,g25800,g14511,g27330,g27393,g26099,g28427,g27258,
    g24681,g16653,g29740,g30005,g28230,g22126,g18128,g21927,g26100,g19588,
    g33416,g32370,g29685,g18245,g27132,g34538,g34330,g18626,g15913,g24730,
    g31992,g31773,g18323,g33841,g33254,g18299,g18533,g28547,g33510,I31247,
    g24765,g17699,g18298,g15073,g27161,g30241,g28729,g18775,g24549,g23162,
    g28226,g27825,g21755,g29334,g29148,g16474,g13666,g23755,g14821,g27259,
    g19749,g32047,g27248,g33835,g9968,g21770,g32205,g21981,g22060,g10902,
    g18737,g27087,g13872,g28572,g27829,g12259,g24504,g22226,g32311,g31295,
    g25207,g22513,g29762,g28298,g18232,g34771,g34693,g29964,g16537,g11027,
    g30235,g28723,g25328,g11890,g7499,g24317,g15797,g18697,g27043,g26335,
    g32051,g31506,I17606,g29587,g18261,g21767,g21794,g15094,g21845,g12043,
    g16303,g24002,g19613,g21990,g11003,g18512,g23990,I27524,g33720,g33161,
    g19560,g15832,g29909,g28435,g27602,g31275,g30147,g34515,g34288,g34414,
    g34206,g31746,g30093,g27375,g26206,g31493,g29791,g32350,g21719,g33493,
    I31161,I31162,g24323,g24299,g13778,g13081,g29569,g29028,g21718,g33465,
    I31022,g31237,g29366,g33237,g32152,g18445,g24775,g17594,g29568,g29747,
    g28286,g32396,g33340,g32222,g21832,g18499,g18316,g33684,g33139,g16840,
    g31142,g22055,g18498,g32413,g31121,g19693,g22111,I31047,g21861,g24653,
    g22070,g13998,g31517,g29849,g26345,g28426,g27257,g33517,I31282,g29751,
    g28297,g29807,g28359,I31311,g29772,g28323,g22590,g19274,g16192,g26849,
    g29974,g29173,g15711,g18611,g15090,g27459,g21926,g15147,g18722,g26399,
    g15572,g25414,g25991,g23389,g29639,g28510,g15109,g26848,I16646,g12413,
    g12343,g26398,g20784,g18432,I24705,g29638,I31051,g21701,I31072,g18271,
    g30082,g29181,g34114,g15108,g21777,g34758,g26652,g10799,g31130,g12191,
    g22067,g22094,g34082,g33709,g30107,g28560,g21251,g13969,I24679,g33362,
    g32259,g11449,g27545,g16483,g18753,g15148,g18461,g31523,g32020,g18342,
    g33523,I31312,g29841,g28371,g19914,g29992,g29012,g34744,g18145,g29510,
    g28856,g32046,g10925,g18199,g22019,g27598,g18650,g18736,g27086,g25836,
    g31475,g29756,g29579,g28457,g17150,I24030,g33475,g16536,g18198,g15059,
    g22018,g15157,g18529,g21997,g32113,g7684,g33727,g33115,g24499,g22217,
    g29578,g33863,g33273,g19594,g11913,g29835,g34141,g16702,g24316,g31222,
    g32282,g31258,g15796,g18330,g32302,g31279,g18393,g24498,g14036,g29586,
    g13821,g12817,g21766,g26833,g26049,g30263,g28773,g32105,g28658,g27563,
    g18764,g16291,g18365,g27158,g26609,g21871,g25107,g17643,g21288,g15840,
    g18132,g26048,g28339,g30135,g28592,g24722,g17618,g34135,I18782,g29615,
    g16673,g18161,g34962,g19637,g26613,g18709,g22001,g22077,g25848,g25539,
    g14190,g27336,g30049,g13114,g18259,g15068,g29746,g28279,g34500,g18225,
    g33351,g32236,g33372,g32285,g18708,g28197,g27647,g25804,g8069,g18471,
    g33821,g33238,g26273,g30048,g29193,g18258,g16634,g16282,g23451,g13805,
    g24199,g24650,g22641,g23220,g24887,I24054,g30004,g28521,I31046,g22624,
    g19344,g21911,g30221,g28700,g31790,g33264,g31965,g31516,g29848,g24198,
    g33790,g33108,g33516,I31276,I31277,g29806,g28358,g29684,g18244,g26234,
    g22102,g24843,I24015,g33873,g33291,g24330,g22157,g24393,g25962,g9258,
    I17552,g24764,g17570,g29517,I31357,g21776,g21785,I27519,g18602,g18810,
    g15757,g18657,g22066,g18774,g18375,g31209,g33422,g32375,g34106,g32248,
    g21754,I27518,g10625,g27309,g26603,g23754,g14816,g28714,g27591,g10699,
    g25833,g14126,I17542,g27288,g26515,g28315,g27232,g33834,g33095,g31208,
    g30262,g32204,g21859,g21825,g21950,g26514,g18337,g28202,g27659,g30033,
    g29189,g28257,g27179,g21858,g29362,g27379,g18171,g30234,g28721,g7450,
    g24709,g16690,g26025,g29523,g28930,g23151,g18994,g28111,g27343,g14296,
    g21996,g24225,g15673,g18792,g15847,g23996,g19596,g24708,g14644,g10610,
    g10605,g16592,g21844,g21394,g13335,g32356,g29475,g14033,g18459,g18425,
    g33905,g33089,g33073,g32386,g25106,g17391,g26541,g34514,g34286,g15851,
    g15872,g18458,g19139,g27374,g33530,g21420,g34507,g34280,g31122,g12144,
    g32182,g31753,g20069,g16312,g33122,g8530,I31027,I24524,g33464,I31016,
    I31017,I16129,g11443,g11411,g20602,g10803,g28150,g12591,g11185,g18545,
    g25951,g24500,g26325,g12644,g24602,g16507,g25972,g18444,g25033,g17500,
    g25371,g24657,g22644,g24774,g16731,g26829,g27669,g17480,g14433,g19333,
    g29347,g29176,g18599,g22307,g20027,g22076,g22085,g26358,g19522,I27349,
    g23025,g16021,g27260,g26766,g32331,g31322,g31292,g29735,g26828,g24919,
    g27668,g23540,g16866,g22054,g28695,g27580,g31153,g12336,g27392,g29600,
    g26121,g20171,g16479,g34541,g34331,g14343,g33409,g32359,I24616,g29952,
    g23576,g27559,g29351,g27525,g27488,g18817,g15912,g14581,g12587,g12428,
    g12357,g18322,g33408,g32358,I31081,g24967,g23197,g10707,g18159,g27558,
    g25507,g18125,g15053,g18532,g26291,g30920,g29889,I24704,g19585,g17180,
    g14202,g16929,g18158,g14257,g21957,g18783,g23957,g29516,g28895,g14496,
    g12411,g12244,g12197,g21739,I31356,g25163,g20217,g18561,g18656,g15120,
    g30121,g28577,g25012,g20644,g18353,g18295,g21738,g17156,g17655,g7897,
    g18680,g15128,g18144,g18823,g34344,g34107,g21699,g28706,g27584,g28597,
    g27515,g18336,g24545,g33474,g28256,g15820,g28689,g27575,g32149,g27042,
    g25774,g30173,g28118,g34291,g34055,g27255,g25936,g28280,g23761,g22131,
    g29834,g28368,g33327,g32208,g34173,g33679,g29208,I27538,I27539,g25788,
    g8010,g32148,g28624,g22357,g28300,g27771,g27270,g32097,g25960,g27678,
    g18631,g32104,g7520,g18364,g32343,g31473,g31283,g30156,g27460,g27686,
    g25946,g24496,g31492,g29790,g24817,g30029,g29164,g33492,g19674,g24322,
    g12939,g27030,g26343,g20977,g10123,g13299,g24532,g22331,g32369,g27267,
    g27294,g9975,g29614,g28860,g30028,g29069,g24977,g23209,g34506,g16803,
    g31750,g30103,g29607,g28509,g18289,I31026,g29320,g29068,g33381,g29073,
    g12065,g18309,g29530,g24656,g29593,g28470,g33091,g32392,g18288,g18224,
    g21715,g22039,g29346,g25173,g12234,g24295,g18571,g18308,g24680,g27219,
    g32412,g24144,g33796,g33117,g19692,g12066,I24555,g29565,g26604,g13248,
    g17469,g13737,g22038,g23551,g10793,g23572,g10917,g12219,g27218,g30927,
    g29910,g18495,g33840,g33253,g29641,g28520,g29797,g28347,g16662,g13697,
    g11166,g28660,g27824,g18816,g32011,g27160,g14163,g10706,g15113,g19207,
    g7803,g18687,g28456,g27290,g17601,g14572,g22143,g19568,g21784,g22937,
    g26845,g24391,g14256,g21956,g18752,g15146,g27455,g26395,g22547,g30604,
    g33522,g18374,g29635,g28910,g21889,g23103,g27617,g26264,g15105,g21980,
    g10624,g28550,g18643,g7469,g32310,g27577,g16204,g27552,g21888,g21824,
    g26633,g34563,g34372,g27201,g26359,g33483,I31112,g26719,g10709,g24289,
    g18669,g32112,g25927,g25004,g32050,g24309,g33862,g33272,g18260,g28243,
    g27879,g24288,g27595,g24224,g18668,g27467,g31949,g18392,g29891,g28420,
    g24308,g21931,g18195,g22015,g18489,g34395,g34193,g31948,g30670,g32096,
    g28269,g27205,g29575,g15881,g18559,g12856,g25491,g23615,g18525,g18488,
    g18424,g28341,g27240,g29711,g33904,g33321,g24495,g28268,g31252,g29643,
    g29327,g29070,g26861,g25021,g25003,g33252,g32155,g13080,g18558,g28655,
    g27561,g30191,g28647,g16233,g29537,g28976,g34191,g16672,g27822,g26389,
    g19949,g18893,g16215,g25981,g24687,g27266,g26612,g26388,g19595,g18544,
    g26324,g32428,g31133,g29606,g28480,g16306,g18713,g13461,g22084,g31183,
    g30249,g26251,g22110,g15167,g24643,g22636,g26272,g33847,g33260,g21860,
    g16513,g13708,g28694,g27579,g29750,g28296,g29982,g23656,g29381,g28135,
    g18610,g15088,g34861,g30247,g28735,g18705,g13887,g25990,g9461,g23497,
    g20169,g33509,I31241,g24669,g22653,g31933,g30926,g29903,g30045,g29200,
    g18255,g18189,g27588,g26690,g15779,g13909,g18679,g31508,g29813,g34389,
    g34170,g13105,g34045,g30612,g26338,g33508,g24668,g21700,g30099,g28549,
    g33872,g33282,g18270,g29796,g28345,g17179,g24392,g22685,g11891,g18188,
    g18124,g21987,g18678,g10802,g16026,g28557,g27772,g34324,g14064,g15081,
    g13393,g16212,g24195,g28210,g32317,g27119,g25877,g30098,g28548,g34701,
    g10721,g20559,g30251,g28745,g34534,g34321,g23658,g14687,g30272,g28814,
    g19206,g15786,g13940,g18460,g18686,g24559,g22993,g18383,g29840,g24488,
    g24016,g14528,g27118,g21186,g11960,g32129,g21943,g25832,g21296,g7879,
    g24558,g22516,g18267,g18294,g15072,g27616,g26349,g26871,g25038,g25020,
    g17654,g32128,I17575,g27313,g29192,g30032,g29072,g21969,g26360,g10589,
    g25573,g30140,g28600,g27276,g9750,g27285,g9912,g29522,g28923,g32323,g31311,
    g24865,g11323,g29663,g34140,g22762,g15651,g21968,g10655,g15672,g27305,
    g10041,g25926,g25005,g24713,g25045,g17525,g18219,g27254,g25935,g30061,
    g33311,g31942,g21855,g34061,g14180,g23855,g22216,g13660,g18218,g21870,
    g28601,g27506,g28677,g27571,g27036,g26329,g29553,g26629,g27177,g27560,
    g26299,g34871,g24189,g31756,g30114,g24679,g13289,g11244,g29949,g23575,
    g32232,g31241,g20188,g18160,g29326,g29105,g28143,g27344,g31780,g30163,
    g25462,I24585,g24188,g22117,g29536,g28969,g22000,g21867,g18455,g24686,
    g24939,g23771,g29757,g28305,I31317,g33350,g32235,g32261,g31251,g18617,
    g18470,g20093,g15372,g33820,g33075,g29621,I24576,g10619,g21714,g23581,
    g20183,g24294,g31152,g25061,g17586,I31002,g18201,g15061,g33846,g33259,
    g21707,g21819,g29564,g18277,g14210,g21910,g26147,g30220,g28699,g28666,
    g27567,g33731,g33116,g28217,g27733,g22123,g21818,I18740,g21979,g16896,
    g27665,g26872,g30246,g28734,g25871,g16281,g18595,g28478,g27007,g18467,
    g18494,g19500,g24219,g26858,g21978,g11967,g18623,g20218,g30071,g29184,
    g17123,g24218,g21986,g34071,g18782,g27485,g28556,g27431,g29509,g32316,
    g31307,g33405,g32354,g21741,g15086,g26844,g25261,g18419,g27454,g26394,
    g22530,g18352,g29634,g29851,g29872,g28401,g28223,g27338,g15104,g34754,
    g18155,g15056,g21067,g18418,g18822,g16713,g32056,g27271,g18266,g11010,
    g8933,g34859,g18170,g10677,g22992,g34370,g34067,g21801,g28110,g27974,
    g21735,g21877,g23801,g34858,g30151,g28607,g30172,g28625,g24915,g23087,
    I31261,g27594,g26721,g28531,g27722,g14378,g22835,g15803,g28178,g27019,
    g18167,g18194,g18589,g22014,g7404,g31787,g34394,g34190,g25071,g33113,
    g31964,g33787,g33103,g32342,g29574,g31282,g30130,g22007,g15850,g29205,
    I27523,g18588,g18524,g28676,g27570,g32145,g14791,g32031,g31372,g24467,
    g13761,g27519,g33357,g32247,g27185,g26190,g25147,g20202,g32199,g30916,
    g18401,g28654,g33105,g26298,g14168,g18477,g26203,g33743,g33119,g16802,
    g18119,g27518,g27154,g9535,g32198,g22116,g16730,g24984,g18118,g21866,
    g21917,g30227,g28708,g31769,g30141,g23917,g33640,g33387,g32330,g31320,
    g29592,g28469,g30059,g28106,g22720,I31316,g30025,g28492,g25151,g16765,
    g15716,g18749,g22041,g26301,g13656,g11144,g18616,g18313,g33803,g33231,
    g24822,g26120,g30058,g29180,g13867,I14198,g18748,g8643,g25367,g21706,
    g18276,g18285,g29350,g26146,g30203,g28668,g18704,g34203,g18305,g33881,
    g33292,g30044,g29174,g18254,g18809,g21923,g22340,g19605,g32161,g22035,
    g28587,g27487,g26290,g18466,g23280,g27215,g27501,g15112,I31271,g30281,
    g28850,g18808,g25420,g24194,g24589,g34281,g34043,g29731,g22142,g27439,
    g34301,g34064,g18177,g18560,g30120,g28576,g28543,g27735,g24588,g32087,
    g34120,g33930,I31342,g32258,g28117,g18642,g15097,g25059,g20870,g33890,
    g33310,g19788,I31031,g16128,g14333,g34146,g33788,g34738,g33249,g32144,
    g34562,g34369,g28569,g27453,g21066,g25058,g23276,g16245,g14278,g32043,
    g31482,g33482,I31106,I31107,g32244,g33248,g32131,g10676,g18733,g15141,
    g27083,g25819,g27348,g33710,g14037,g22130,g27284,g9908,g24864,g11201,
    g22193,g19880,g28242,g27769,g21876,g21885,g26547,g13283,g10654,g11023,
    g15857,g23885,g27304,g24749,g17511,g32069,g10878,g12284,g14654,g24313,
    g22165,g15594,g18630,g21854,g15793,g18693,g23854,g31778,g24748,g17656,
    g32068,g31515,g33081,g32388,g17193,g21763,g18166,g24285,g25902,g24398,
    g18665,g31786,g30189,g25957,g17190,g24704,g17593,g25377,g33786,g33130,
    g24305,g16737,g26572,g22006,g28639,g27767,g24900,I24067,g33647,g33390,
    g32337,g31465,g27139,g28293,g33356,g32245,g22863,g27653,g28638,g27551,
    g32171,g31706,g18476,g18485,g29787,g28334,g26127,g27138,g28265,g34661,
    g18555,g18454,g25290,g14216,g21916,g30226,g28707,g18570,g18712,g33233,
    g32094,g31182,g30240,g27333,g24642,g34226,g33914,g14587,g10584,g10567,
    g29743,g28206,g34715,g34481,g34404,g32425,g31668,g26103,g34572,g10543,
    g8238,g26095,g11923,g27963,g25952,g29640,g28498,g25366,g29769,g28319,
    g18239,g21721,g33331,g32216,g27664,g18567,g18594,g12858,g31513,g32010,
    g31785,g33513,I31262,g29803,g28414,g18238,g26181,g26671,g28586,g27484,
    g24630,g23255,g31961,g31751,g33897,g33315,I18785,g31505,g28442,g27278,
    g33505,I31221,g18382,g24009,g19671,g33404,g32353,g29881,g21773,g18519,
    g11016,g8984,g21942,g13525,g18176,g18185,g22063,g18675,g34385,g34168,
    g33717,g14092,g24008,g32086,g30095,g28545,g31212,g28116,g27366,g18518,
    g18154,g27312,g12019,g24892,g11559,g24476,g18879,I31337,g16611,g27115,
    g11893,g13830,g11543,g11424,g11395,g22873,g19854,g25551,g23822,g18637,
    g25572,I24699,I24700,I31171,g30181,g28636,g30671,g29319,g32322,g31308,
    g24555,g23184,g29662,g9217,g21734,g32159,g24712,g29890,g28419,g24914,g8721,
    g21839,g21930,g25127,g13997,g21993,g32158,g22209,g19907,g15856,g10666,
    g33723,g14091,g28237,g21838,g22834,g15880,g31149,g29508,g21965,g15149,
    g26088,g26024,g22208,g19906,g29710,g28035,I26530,I26531,g29552,g33433,
    g32238,g23131,g13919,g32295,g27931,g10841,g29204,g31148,g30190,g28646,
    g13042,g16199,g25103,g27184,g26628,g16736,g18501,g12854,g18729,g15139,
    g22021,g27674,g26873,g25980,g18577,g33104,g26296,g25095,g23319,g33811,
    g33439,g33646,g33389,g19767,g16810,g32336,g34520,g34294,g23619,g19453,
    g33343,g32227,g21557,g12980,g18728,g18439,g30089,g28538,g24941,g23171,
    g26126,g30211,g28685,g11939,g23618,g19388,g25181,g23405,g16843,g18438,
    g34211,g33891,g26250,g13383,g24675,g17568,g29647,g28934,g30024,g28497,
    g33369,g32277,g17726,g16764,g13030,g22073,g18349,g14586,g11953,g11970,
    g13294,g29380,g28134,g33368,g32275,g34860,g16869,g27692,g26392,g28130,
    g27353,g28193,g26339,g25931,g24574,g18906,g13568,g18348,g24637,g16586,
    g19521,g22122,g12761,g18284,g15071,g16868,g34497,g28165,g28523,g27704,
    g18304,g29182,g29651,g33412,g32362,I31322,g16161,g15611,g15722,g18622,
    g22034,g15080,g12855,g18566,g30126,g28582,g14615,g10604,g10587,g27214,
    g34700,g34535,g31229,g30288,g10720,g21815,g30250,g28744,g27329,g12052,
    g32309,g27207,g33896,g33314,g31228,g27539,g29331,g29143,g32224,g34658,
    g23187,g13989,g26855,g21975,g27328,g12482,g25089,g23317,g32308,g31293,
    g20215,g29513,g28448,g18139,g27538,g18653,g24501,g14000,g24729,g25088,
    g13093,g11160,g17153,I24033,g18138,g21937,g34338,g34099,g24728,I17585,
    I31336,g15650,g34969,g10684,g28703,g27925,g18636,g18415,g31310,g30157,
    g18333,g30060,g29146,g21791,g28253,g23719,g21884,g11915,g34968,g23884,
    g30197,g28661,g31959,g33379,g19462,g7850,g14182,g14177,g25126,g16839,
    g25987,g13277,g28236,g34870,g34527,g34303,g24284,g18664,g27235,g25910,
    g24304,g26819,g27683,g25770,g24622,g19856,g33742,g26257,g31944,g31745,
    g11037,g18576,g18585,g14193,g18484,g22109,g32260,g31250,g28264,g34503,
    g34278,g34867,g34826,g25969,g9310,g18554,g29620,g33681,g33129,g22108,
    g18609,g32195,g30734,g24139,g25968,g25215,g18312,g33802,g33097,g33429,
    g32231,g33857,g33267,g29646,g30315,g22864,g18608,g15087,g27407,g18115,
    I27534,g33730,g32016,g33428,g32230,g34707,g30202,g28667,g25870,g24840,
    g30257,g28750,g25411,I24546,g26094,g31765,g30128,g24415,g7763,g24333,
    g29369,g28209,g14222,g21922,g22982,g19535,g30111,g28565,g18745,g33690,
    g33146,g30070,g29167,g34111,g33733,g18799,g22091,g23531,g10760,g13853,
    g18813,g30590,g21740,g16599,g26019,g25503,g18798,g28542,g27405,g31504,
    g29370,g28453,g27582,g27206,g33504,g24664,g22652,g29850,g28340,g19911,
    g14707,g34741,g16598,g15810,g13524,g17091,g18184,g21953,g18805,g18674,
    g23373,g13699,g30094,g28544,g25581,g25450,g32042,g27244,g21800,g16288,
    g23208,g29896,g27114,g32255,g31248,g31129,g32189,g30824,g21936,g18732,
    g27435,g18934,g24554,g22490,g27107,g32270,g31254,g16125,g16532,g25818,
    g8124,g28530,g27383,g31128,g12187,g32188,g27586,g25979,g24517,g28346,
    g27243,g7251,g24312,g18692,g18761,g33245,g32125,g24608,g25978,g9391,g13313,
    g15967,g30196,g28659,g31323,g30150,g29582,g27766,g31299,g30123,g17192,
    g34196,g21762,g21964,g25986,g32030,g24921,g23721,g31298,g30169,g34526,
    g34300,g18400,g10873,g26077,g24745,g29627,g28493,g18214,g28292,g23781,
    g29959,g28953,g22862,g27031,g18329,g25067,g25094,g23318,g18207,g26689,
    g15754,g29378,g13808,g18539,g11036,g26280,g18328,g27263,g25940,g21909,
    g31232,g30294,g25150,g22040,g25801,g26300,g34866,g34819,g28136,g27382,
    g18538,g27332,g12538,g29603,g24674,g29742,g28288,g21908,g33697,g33160,
    g30001,g28490,g31995,g33856,g33266,g26102,g12135,g31261,g14754,g26157,
    g27406,g27962,g25954,g27361,g33880,g33290,g18241,g34706,g34496,g21747,
    g32160,g31001,g30256,g28749,g25526,g23720,g28164,g26231,g33512,g14913,
    g27500,g29857,g28386,g15817,g14614,g11975,g11997,g24761,g22751,g21814,
    g18771,g16023,g14583,I14225,g18235,g21751,g21807,g21772,g26854,g15783,
    g21974,g22062,g18683,g25866,g24400,g27221,g28327,g27365,g29549,g34102,
    g26511,g19265,g34157,g33794,g10565,g8182,g28537,g31499,g29801,g33499,
    I31191,g14565,g11934,g11952,g29548,g24329,g30066,g28518,g22851,g28108,
    g30231,g28718,g15823,g34066,g10034,g25077,g23297,g33498,g23265,g24328,
    g28283,g18515,g23416,g20082,g18414,g31989,g31770,g14641,g11994,g12020,
    g28303,g27106,g21841,g21992,g34876,g18407,g25923,g24443,g31988,g31768,
    g33722,g33175,g33924,g32419,g15966,g28982,g31271,g29706,g12812,g34763,
    g15631,g27033,g25767,g27371,g32418,g31126,g26287,g27234,g25102,g21835,
    g32170,g31671,g13567,g22047,g26307,g26085,g11906,g29626,g28584,g33461,
    g16669,g33342,g32226,g29323,g23007,g31145,g18441,g18584,g24771,g18206,
    g29533,g28958,g12795,g16668,g16842,g14546,g33887,g33298,g18759,g22051,
    g22072,g18725,g32167,g32194,g25876,g33529,I31201,g27507,g18114,g28192,
    g18758,g26341,g24746,g18435,g33528,g11370,g19661,g33843,g33256,g21720,
    g33330,g32211,g26156,g18107,g28663,g27566,g32401,g31116,g34076,g33694,
    g30596,g30279,g26180,g26670,g21746,g33365,g32267,g32119,g30243,g28731,
    g31132,g29504,g18744,g34054,g31960,g31749,g33869,g33279,g14537,g10550,
    g10529,g18345,g19715,g29856,g28385,g21465,g16155,g18399,g29880,g33868,
    g33278,g26839,g27541,g26278,g30269,g28778,g22846,g21983,g28553,g25456,
    I24579,g18398,g29512,g32313,g31303,g21806,g26838,g18141,g30268,g28777,
    g18652,g18804,g15163,g34341,g34101,g25916,g24432,g16610,g16705,g17152,
    g31225,g30276,g32276,g34655,g27359,g30180,g28635,g27325,g12478,g29359,
    g31471,g29754,g32305,g31287,g32053,g14176,g33471,I31052,g34180,g33087,
    g32391,g18263,g32254,g31247,g27535,g26487,g15702,g27434,g27358,g25076,
    g25085,g18332,g19784,g28252,g27159,g12920,g18135,g8461,g25054,g24725,
    g19587,g30930,g29915,g32036,g31469,g27121,g29316,g28528,g19354,g33244,
    g32177,g30608,g18406,g13349,g11780,I31167,g26279,g18361,g24758,g23130,
    g34667,g34694,g17405,g13137,g34965,g30131,g28589,g31069,g29793,g29989,
    g29006,g18500,g22020,g27682,g25777,g23165,g13954,g28183,g27024,g28673,
    g33810,g33427,g27291,g11969,g29611,g28540,g33657,g26286,g29988,g29187,
    g29924,g13031,g34487,g34416,g13566,g22046,g26306,g24849,g33879,g33289,
    g24940,g24399,g26363,g30210,g28684,g34557,g34352,g23006,g19575,g23475,
    g19070,g33878,g33288,g18221,g22113,g21863,g26815,g24141,g34279,g34231,
    g11139,g33886,g33297,g27134,g30278,g28818,g27029,g26327,g18613,g31792,
    g30214,g32166,g31007,g32009,g31782,g25993,g31967,g31755,g31994,g31775,
    g22105,g27028,g26342,g32008,g31781,g25965,g29650,g28949,g29736,g28522,
    g16160,g29887,g28417,g21703,g24332,g18106,g20135,g16258,g18605,g13415,
    g21347,g13333,g11755,g33425,g32380,g28213,g27720,g15679,g18812,g18463,
    g33919,g33438,g24406,g13623,g29528,g24962,g23194,g29843,g28373,g21781,
    g29330,g29114,g16617,g25502,g15678,g18951,g30187,g28643,g18371,g28205,
    g27516,g18234,g34187,g17769,g21952,g28311,g23372,g16448,g29869,g21821,
    g17768,g13325,g18795,g29868,g27649,g10820,g34143,g16595,g21790,g24004,
    g33086,g32390,g27648,g24221,g27491,g26486,g18514,g29709,g21873,g18507,
    g22027,g23873,g15875,g30168,g28623,g29708,g33817,g33235,g11115,g33322,
    g32202,g34410,g34204,g27981,g26751,g25815,g31125,g29502,g32176,I31166,
    g26223,g31977,g31764,g33532,g33901,g33317,g34479,g34403,g34666,g25187,
    g12296,g18163,g15837,g32154,g31277,g34363,g34148,g25975,g34217,g22710,
    g19358,g30015,g29040,g21834,g22003,g34478,g34402,g28152,g26297,g26084,
    g28846,g24812,g19855,g33353,g32240,g25143,g34486,g34412,g18541,g33680,
    g33128,g18473,g27262,g26179,g12794,I17529,g34556,g34350,g18789,g21453,
    g22081,g29602,g29810,g28259,g29774,g28287,g29539,g26178,g27633,g13076,
    g21913,g29375,g13946,g30223,g28702,g11489,g11394,g11356,g18788,g18724,
    g25884,g11153,g18359,g34223,g18325,g26186,g24580,g18535,g18434,g18358,
    g31966,g31754,g30084,g28534,g27521,g29337,g29166,g17786,g30110,g28564,
    g25479,g34084,g15075,g12850,g31017,g29479,g34110,g33732,g25217,g12418,
    g33364,g32264,g18121,g22090,g30179,g28634,g24507,g22304,g18344,g19581,
    g15843,g34179,g21464,g16181,g28020,g28583,g30178,g28632,g9479,g24421,
    g34178,g34740,g16616,g10756,g18682,g30186,g28641,g27247,g18291,g24012,
    g17182,g21797,g34186,g34685,g14164,g25580,g18173,g27389,g34953,g27045,
    g31309,g30132,g32083,g32348,g23292,g19879,g25223,g22523,g16704,g27612,
    g25887,g31224,g30280,g32284,g31260,g28113,g26423,g19488,g27099,g14094,
    g15822,g27388,g27324,g32304,g31284,g30936,g28282,g23762,g12099,g27534,
    g27098,g25868,g28302,g23809,g25084,g27251,g27272,g25110,g16808,g19384,
    g18760,g18134,g25922,g24959,g34334,g34090,g24788,g11384,g31495,g24724,
    g17624,g29599,g33495,g22717,g16177,g24325,g25179,g16928,g26543,g12910,
    I27503,g18506,g22026,g27462,g33816,g33234,g29598,g28823,g16642,g25178,
    g20241,g15589,g32139,g27032,g34964,g33687,g33132,g31976,g31762,g31985,
    g19735,g27140,g25885,g30216,g28691,g27997,g26813,g28768,g15836,g31752,
    g30104,g34216,g31374,g29748,g29322,g33374,g32289,g16733,I18671,g29532,
    g29901,g28429,g32333,g31326,g15119,g16238,g11441,g11355,g11302,g25417,
    g23474,g24682,g22662,g22149,g29783,g28329,g21711,g26123,g15118,g34909,
    g34856,g24291,g30000,g23685,g29656,g28515,g34117,g15749,g18649,g22097,
    g27360,g33842,g33255,g18240,g15066,g22104,g17149,g33392,g32344,g18648,
    g18491,g31489,g26230,g25964,g33489,I31141,g21606,g15959,g27162,g34568,
    g34379,g34747,g23606,g16927,g29336,g15704,g30242,g28730,g18604,g21303,
    g16485,g18755,g31525,g29892,g31488,g31016,g29478,g33525,g33488,g28249,
    g27152,g15809,g18770,g15153,g20783,g18563,g18981,g11206,g21750,g28248,
    g27150,g29966,g23617,g28710,g27589,g15808,g21982,g27451,g26391,g19593,
    I26948,g23381,g27220,g33830,g29631,g32312,g31302,g32200,g27468,g33893,
    g33313,g28204,g26098,g27628,g34751,g29364,g27400,g10827,g25909,g32115,
    g25543,g23795,g12220,g27246,g33865,g33275,g21796,g30230,g28717,g25908,
    g24782,g18767,g15150,g18794,g34230,g18395,g12849,g32052,g31507,g18262,
    g22133,g25569,I24685,g21840,g15099,g25568,g18633,g17133,g34841,g34761,
    g18191,g18719,g22011,g15154,g15874,g24649,g29571,g28452,g11114,g31270,
    g29692,g16519,g16176,g14596,g16185,g25123,g18718,g15693,g18521,g31188,
    g25814,g24760,g27370,g31124,g32184,g30611,g17424,g33124,g24903,g28233,
    g27827,g16518,g28182,g25772,g24944,g24934,g28672,g24755,g16022,g27151,
    g24578,g16637,g22310,g18440,g13345,g11773,g26275,g30007,g29141,g11025,
    g18573,g29687,g22112,g18247,g29985,g21862,g22050,g23553,g19413,g18389,
    g29752,g28516,g29954,g21949,g15712,g18612,g15914,g25992,g18388,g19660,
    g12001,g18324,g24794,g11414,g31219,g30265,g34116,g33933,g24395,g25510,
    I24619,g18701,g26684,g25407,g21948,g22096,g32400,g18777,g18534,g32013,
    g30041,g28511,g18251,g21702,g31218,g30271,g16729,g18272,g21757,g25579,
    g30275,g28816,g27227,g33837,g33251,g32207,g31221,g26517,g15708,g34746,
    g34493,g34273,g25578,g15567,g27025,g26334,g24191,g24719,g18462,g25014,
    g17474,g32328,g29668,g28527,g29842,g28372,g27540,g23564,g16882,g27058,
    g30035,g22539,g18140,g34340,g34100,g27203,g26130,g24890,g29525,g21847,
    g34684,g14178,g13833,I18819,g26362,g19557,g27044,g31470,g29753,g23397,
    g11154,g33470,g33915,g33140,g32241,g31244,g26165,g11980,g10998,g18766,
    g13048,g23062,g27281,g9830,g24861,g24573,g17198,g34517,g34290,g28148,
    g27355,g14233,g21933,g27301,g11992,g27957,g25947,g7804,g25041,g23261,
    g13221,g27120,g25878,g29865,g21851,g21872,g23872,g15883,g18360,g31467,
    g30162,g31494,g29792,g28343,g27380,g19655,g33467,I31032,g33494,g24324,
    g27146,g27645,g26863,g24974,g24957,g18447,g30193,g28650,g24777,g11345,
    g27699,g26396,g13850,g18162,g25983,g29610,g28483,g30165,g28619,g22129,
    g34523,g22002,g22057,g15159,g17317,g13124,g22128,g33352,g32237,g16636,
    g18629,g25142,g18451,g26347,g18472,g32414,g33418,g32372,g33822,g18220,
    g26253,g30006,g29032,g31266,g30129,g21452,g18628,g15095,g27427,g27450,
    g17057,g24140,g22299,g19999,g29686,g18246,g21912,g29383,g28138,g30222,
    g28701,g34863,g28133,g27367,g22298,g19997,g28229,g27345,g19487,g29938,
    g23552,g26351,g28228,g27126,g25130,g23358,g26821,g24821,g27661,g27547,
    g18591,g31167,g18776,g18785,g21756,g18147,g25165,g14062,g30253,g28746,
    g16484,g18754,g31524,g33524,g18355,g33836,g33096,g21780,g29875,g28403,
    g32206,g30609,g26516,g13507,g27481,g30600,g30287,g18825,g18950,g11193,
    g18370,g31477,g29763,g33401,g32349,g33477,I31082,g20162,g8737,g30236,
    g28724,g14148,g29837,g28369,g14097,g21820,g11163,g9906,g18151,g31118,
    g29490,g18172,g15058,g28627,g27543,g32114,g30175,g28629,g32082,g33864,
    g33274,g27127,g21846,g28112,g27352,g32107,g15653,g24629,g23396,g20051,
    g18367,g18394,g31313,g30160,g24451,g21731,g24220,g20628,g27490,g13541,
    g30264,g28774,g34063,g13473,g30137,g28594,g19601,g16198,g24628,g32345,
    g34137,g31285,g30134,g34516,g34289,g27376,g27385,g29617,g31305,g29741,
    g27103,g33305,g31935,g22831,g19441,g23691,g14731,g26542,g13102,g34873,
    g26021,g18420,g15852,g13820,g27095,g18319,g33809,g33432,g33900,g33316,
    g33466,g16184,g16805,g21405,g13377,g16674,g29201,g32141,g22316,g18318,
    g18446,g33808,g33109,g24785,g18227,g7777,g27181,g30209,g28682,g21334,
    g33101,g32398,g19791,g14253,g24754,g19604,g29595,g28475,g29494,g30208,
    g28681,g16732,g21929,g32263,g18540,g10896,g22056,g26274,g29623,g28496,
    g32332,g31325,g21928,g22080,g25063,g13078,g24858,g29782,g28328,g18203,
    g26122,g24557,g16761,g29984,g34542,g34332,g21187,g12931,g29352,g25873,
    g24854,g18281,g27520,g21787,g15091,g15115,g21287,g18301,g30607,g30291,
    g32049,g26292,g33693,g33145,g18377,g19556,g11932,g30073,g22145,g18120,
    g26153,g24565,g18739,g21302,g22031,g27546,g30274,g28815,g31166,g34073,
    g16207,g27211,g32048,g31498,g21743,g21827,g11029,g17753,g13281,g18146,
    g18738,g15142,g13029,g8359,g15745,g18645,g15100,g30122,g28578,g24420,
    g23997,g24319,g29853,g16538,g17145,g26635,g25321,g11028,g18699,g34565,
    g34374,g15813,g31485,g29776,g29589,g33892,g33312,g18290,g17199,g24318,
    g33476,g33485,I31121,g21769,g30034,g29077,g22843,g24227,g18698,g15131,
    g25453,g29588,g29524,g29836,g28425,g21768,g21803,g28245,g15805,g28626,
    g27542,g30153,g28610,g28299,g22132,g29477,g14090,g32273,g31255,g32106,
    g18427,g14681,g19740,g20203,g18366,g21881,g27658,g22491,g18632,g25905,
    g24879,g17365,g33074,g32387,g34136,g33239,g32117,g25530,g23750,g27339,
    g29749,g28295,g29616,g7511,g26711,g25446,g31238,g29583,g32234,g25122,
    g23374,g18403,g18547,g25565,g13013,g24301,g28232,g27732,g16259,g13491,
    g22087,g30164,g28618,g31941,g33941,g33380,g18226,g15064,g21890,g13604,
    g31519,g29864,g18715,g27968,g25958,g28697,g27581,g31185,g18481,g33519,
    I31291,g29809,g28362,g24645,g22639,g28261,g27878,g26606,g28880,g18551,
    g22043,g26303,g31518,g18572,g33518,g29808,g28361,g21710,g24290,g29036,
    g27411,g20083,g24698,g22664,g21779,g26750,g24514,g12527,g23779,g18127,
    g22069,g25408,g30109,g28562,g26381,g34109,g29642,g27954,g33883,g33294,
    g21778,g22068,g26091,g18490,g30108,g28561,g32163,g32012,g24427,g21786,
    g27503,g30283,g28851,g18784,g15155,g18376,g18385,g29733,g18297,g17810,
    g18103,g10626,g34492,g13633,g25164,g16883,g21945,g28499,g27982,g18354,
    g29874,g28402,g21826,g21999,g26390,g31501,g18824,g27315,g12022,g33501,
    g29630,g28212,g24403,g29693,g28207,g30982,g34750,g16759,g18181,g21998,
    g18671,g34381,g34166,g23998,g27202,g30091,g32325,g31316,g29665,g16758,
    g24226,g13832,g28722,g27955,g30174,g28628,g29008,g12979,g24551,g17148,
    g24572,g33349,g32233,g25108,g23345,g21932,g32121,g18426,g33906,g33084,
    g13247,g29555,g29004,g21513,g16196,g18190,g22010,g23513,g19430,g34390,
    g34172,g10856,g11045,g15882,g27384,g29570,g29712,g33304,g32427,g14261,
    g18520,g21961,g22079,g27094,g30192,g28649,g13324,g29907,g32291,g31268,
    g16804,g21404,g28199,g27479,g22078,g23404,g20063,g32173,g18546,g25982,
    g18211,g15062,g21717,g15051,g28198,g26649,g24297,g22086,g25091,g20095,
    g8873,g29567,g29594,g28529,g31139,g12221,g28330,g27238,g26252,g11032,
    g34483,g34406,g18497,g32029,g31318,g24671,g14831,g22125,g28172,g27526,
    g34862,g29519,g32028,g19578,g16183,g33415,g32368,g22158,g13698,g14316,
    g33333,g32218,g18700,g15132,g18126,g15054,g18659,g18625,g15092,g18987,
    g29518,g28906,g18250,g24931,g23153,g15114,g25192,g20276,g26847,g34948,
    g18658,g15121,g27457,g26397,g19475,g15082,g23387,g16506,g31963,g30731,
    g29637,g19530,g7781,g34702,g34537,g15107,g34757,g17783,g25522,g24190,
    g18339,g18943,g29883,g18296,g21811,g28225,g27770,g23104,g23811,g23646,
    g16959,g18644,g15098,g28471,g16221,g18338,g30564,g9967,g28258,g27182,
    g21971,g34564,g34373,g15849,g31484,g29775,g24546,g22447,g33484,g16613,
    g15848,g19275,g7823,g27256,g25937,g19746,g28244,g27926,g34183,g18197,
    g22017,g15652,g15804,g7673,g25949,g24701,g27280,g9825,g31312,g30136,g29577,
    g30062,g13129,g27300,g12370,g10736,g31115,g29487,g18411,g25536,g23770,
    g25040,g34509,g34283,g21850,g28602,g27509,g23412,g28657,g27562,g25904,
    g14001,g19684,g34508,g34282,g10528,g34872,g24700,g24659,g12459,g12306,
    g12245,g26205,g23229,g29349,g22309,g20658,g18503,g22023,g26311,g24658,
    g22645,g22308,g28171,g27016,g33798,g33227,g21716,g30213,g28688,g24296,
    g18581,g18714,g26051,g24896,g18450,g31184,g34213,g18315,g33805,g33232,
    g24644,g29622,g29566,g18707,g15134,g18819,g18910,g16227,g18202,g30047,
    g29109,g18257,g26780,g30205,g28671,g32191,g27593,g18818,g15165,g18496,
    g34205,g31934,g31670,g18111,g21959,g21925,g26350,g25872,g28919,g27663,
    g12369,g28458,g24197,g24855,g16163,g14254,g22752,g15792,g15613,g18590,
    g21958,g21378,g7887,g23050,g28010,g30051,g28513,g26846,g18741,g15143,
    g34072,g23386,g20034,g30592,g30270,g18384,g29636,g21742,g17752,g27480,
    g34756,g28599,g27027,g21944,g33400,g32347,g29852,g14599,g15812,g13319,
    g27314,g12436,g24503,g22225,g27287,g26545,g32045,g31491,g33329,g32210,
    g31207,g30252,g18150,g10657,g18801,g15160,g18735,g25574,g27085,g25835,
    g32324,g31315,g29664,g33328,g32209,g21802,g22489,g12954,g21857,g16535,
    g20581,g10801,g10970,g23857,g13059,g13025,g30152,g28609,g24581,g24714,
    g32098,g24450,g21730,g24315,g21793,g32272,g22525,g13006,g28159,g18196,
    g22016,g28125,g27381,g15795,g28532,g27394,g34396,g34194,g24707,g13295,
    g29361,g29576,g29585,g21765,g27037,g18526,g27269,g25943,g29554,g28997,
    g23690,g14726,g19372,g26020,g33241,g34413,g13176,g11044,g27341,g29609,
    g28482,g27268,g25942,g32032,g31373,g25780,g25532,g25527,g15507,g32140,
    g18402,g18457,g24590,g29608,g28568,g27180,g16097,g20094,g27335,g12087,
    g13738,g25152,g23383,g22042,g26302,g26357,g29799,g28271,g30583,g29355,
    g16760,g27667,g26361,g18706,g25834,g13290,g29798,g28348,g22124,g27131,
    g30046,g29108,g18256,g29973,g28981,g18689,g15129,g31991,g33515,I31272,
    g33882,g33293,g18280,g29805,g28357,g33414,g32367,g22686,g19335,g22939,
    g18688,g18624,g32162,g31002,g18300,g24196,g33407,g32357,g34113,g27502,
    g11427,g22030,g22938,g19782,g27557,g22093,g23533,g19436,g11366,g27210,
    g21298,g29732,g28289,g27734,g21775,g12461,g12415,g13632,g18157,g15057,
    g23775,g14872,g22065,g34743,g28571,g27458,g24402,g29761,g28310,g18231,
    g21737,g32246,g31246,g22219,g19953,g25928,g25022,g8583,g27286,g33441,
    g32251,g31206,g30260,g10656,g27039,g22218,g19951,g28495,g27012,g32071,
    g27236,g21856,g14295,g21995,g31759,g23856,g14680,g12024,g12053,g33759,
    g33123,g24001,g21880,g29329,g25113,g23346,g18511,g29207,g25787,g24792,
    g32147,g18763,g31758,g30115,g33114,g24706,g15910,g26249,g33758,g33133,
    g22160,g27601,g33082,g32389,g21512,g16225,g29328,g27677,g13021,g23810,
    g23786,g29538,g11127,g24923,g23129,g25105,g13973,g10966,g31744,g30092,
    g22681,g22663,g26204,g24624,g16524,g24300,g15123,g26779,g24497,g33345,
    g32229,g32151,g32172,g31940,g18456,g33849,g33262,g30027,g29104,g33399,
    g32346,g21831,g26778,g25501,g34662,g16845,g11956,g18480,I28566,I30330,
    I31859,g16926,I25736,I31858,g24148,g26879,g32455,g33951,g20214,g20199,
    I22298,I31844,g22535,g24018,g26874,I31838,I31839,g11448,g8913,g24609,
    g24965,g23825,g24468,g22400,g14419,g14397,g11999,I18495,g32426,g30613,
    g22540,g14450,g14420,g12025,I18543,g24363,g24478,g22450,g24433,I26643,
    I18492,g14538,g14513,g14446,g7223,g7201,g30317,I28567,g24460,g21384,g21363,
    I22830,g24661,g26052,g8921,I12902,I12903,g24620,g25974,g22585,I30124,
    I12583,g25856,g24591,g22488,g25504,g25141,I18452,g14514,g14448,g14418,
    g9483,g22537,g26657,g26878,g24566,g24678,g9536,I29986,g22522,I31854,g33957,
    I31868,I31869,I24117,g25010,g33956,I31863,I31864,g16876,I18449,g14512,
    g14445,g14415,I30728,I30745,I30746,I28147,g24561,g28220,g20522,g21652,
    g25575,I23163,g29520,g11372,I12611,I30761,I30400,g24880,g25953,g20198,
    g20185,I22280,g26616,I23755,g29496,g24447,g21432,g21416,I22912,I25612,
    I25613,g10821,g8790,I12782,I12783,I30399,g8904,g13091,g28191,g32845,g32780,
    I23162,g20271,g20150,g20134,g10511,I31873,I26644,I30740,I30741,g19525,
    g16811,g26636,g25577,I26741,I26742,I29351,g33953,I31848,I31849,g24544,
    g25996,g11184,g14364,g14337,g11958,I18421,I30760,g25576,g29486,g24547,
    g26053,g14539,g14515,g14449,I30755,g25805,I30262,I30718,g32585,g24652,
    g25995,g24457,g11380,g20184,g20170,I22267,g33952,I31843,g8905,g29529,
    g32520,g24471,g14396,g14365,g11976,I30727,g24444,I23756,g9012,g32910,
    g33958,g22531,g22669,g13914,I30055,I30735,g14416,g14394,g11995,g26866,
    g14187,g8871,g11771,g22514,g14393,g14362,g11972,g28186,g21555,g21364,
    g21357,I30750,I30751,I30054,I30734,g21401,g21385,I22852,I30756,g24145,
    I30469,I30468,g29482,g34912,I30717,g9055,g13938,g11213,g11191,g22517,
    g14447,g14417,g14395,g14334,g14313,g11935,I18385,g24584,g25984,I31874,
    g28031,g27223,g27141,g8956,g21658,I30123,g8957,g21655,g21415,g21402,I22880,
    g22524,I29985,I22958,g21603,g21386,g21365,I26523,I30193,g20371,g20161,
    g20151,I31853,g33955,g21509,g21356,g21351,g25839,g9013,I29352,g25791,
    g29914,g14413,g14391,g14360,g33954,I26522,I30192,g21462,g21433,g29495,
    g32715,g29489,g29488,g13972,g11232,g11203,g8863,g21429,g21338,g21307,
    g32650,g20236,g20133,g20111,g25821,I30331,g13794,g29485,g29501,I18417,
    g14444,g14414,g14392,g13858,g14568,g14540,g14516,g14361,g14335,g11954,
    g21459,g21350,g21339,g10819,I30261,I14817,I14818,g11566,g11435,g12169,
    I22761,I22760,I13443,I13442,I14185,g16719,g13700,I14518,I14516,g17595,
    g14367,g22984,I12346,I12344,I15299,I15300,g17790,g14820,g17761,g14780,
    I14883,g19474,g11426,g11190,g9852,I25908,I25909,I15089,I15087,g22853,
    g21353,I15088,g24916,g19450,g25779,g24362,g12084,g22836,g21330,g20076,
    g13795,g15744,g13119,g15730,g13100,g23132,g19932,I22683,g27796,I13391,
    I13392,I11865,I11866,g15719,g14490,I20165,g16246,g14489,g9694,g20838,
    g23623,g24942,g20039,I26459,g14306,g13256,g14830,g12211,I32431,g34056,
    g34051,I13510,I13511,I20222,g16272,I20221,g12323,g14408,g17312,I25244,
    I25242,g11968,g9334,g13968,g11255,g12716,g7142,I15242,I15243,g24917,g25018,
    g24918,g17284,g13855,g10922,I13110,I13109,g22642,g13870,g13527,I22973,
    I22974,g14317,g17217,g16628,g11207,I23119,I23118,g12000,g22874,g7352,
    g11312,g14686,g12059,I12840,g9640,g16776,g13772,g10715,g11707,I18530,
    I18529,I14609,g8678,I13334,g13257,g27933,g17814,g14854,g17605,g17581,
    g11979,g13496,g11590,g12639,g22712,g23010,I12288,I12289,g24601,g11747,
    g24677,g21388,g17712,g14425,g12416,g11626,g8958,g13067,I18635,g14713,
    I18633,g10617,g16319,I32187,I32185,I12252,I12251,g12553,g10266,g22941,
    I17406,I17404,g10341,g24924,g24905,g12014,g11658,g11527,g10623,g17675,
    g14399,I22800,I22801,I13751,I13749,g12755,g10491,I14400,I14398,g12116,
    g12680,g13866,g11194,I18537,I18536,g13937,g12632,g11715,g11537,I22972,
    g15787,g15781,g15753,g13131,I13390,g11846,I13509,I14734,I14735,g12340,
    g12035,g11692,I15298,I13402,I13403,g20186,g8177,g14379,g17287,g17493,
    I12205,I12203,g10759,g9755,g17492,g13066,g20173,g23379,g11679,g10421,g7227,
    I32186,g13854,I14481,I14482,I14991,g13511,g20216,I20487,I20488,g11933,
    g11951,g9762,g12222,g22852,g11653,g11729,g25002,I29297,g12117,I29295,g8906,
    I26460,I22946,I22944,g14642,I15287,I14206,I14204,g16956,g13824,I26093,
    g13539,I15307,I15306,g23195,g10695,I15241,g13475,g13495,g13057,g13459,
    I15194,I15195,g20011,g23167,I23979,I23980,I15341,I15340,g12604,g12798,
    g21301,g31997,g22306,g30580,g11610,I14399,I13044,I13045,g22921,g15715,
    g14248,g24621,g12700,g12515,g17608,g12067,g12969,I18634,I15335,I15333,
    I31984,I31985,g14570,g13993,I23963,g13631,I23961,I13519,I13520,g21124,
    g17393,I14332,g9966,I14330,g13667,g11119,g12101,g20007,I23585,g13739,
    g21294,g13210,I32757,I32758,g16625,g17732,I15263,I15264,g11279,g14519,
    g11225,I29296,g12317,I25219,g24972,g24950,g24906,I26419,g14247,I26417,
    I22755,I22753,g12073,g11669,g14529,I26418,g12374,g12255,g16296,g13501,
    I24462,I24463,g7133,I11825,I11826,g12464,g12797,I22794,I22792,I22845,
    g12113,I22844,I12204,g30573,g12292,I13140,I13141,g12153,I24364,I24365,
    I22899,g12193,g8829,I22762,g12780,I20205,I20203,I14992,I14993,I22719,
    I22717,g9904,I13444,g7661,I13453,I13452,I22718,g33394,g11169,I14229,I14230,
    I29315,g12154,I29313,I15168,g9823,I15166,g13884,g11410,g20717,I13111,
    I15363,I12402,I12403,g11479,g13479,g12686,g12590,g12526,I12373,I12374,
    I32517,g34424,I32516,g10622,g13478,g12511,g12460,g12414,g12344,I13565,
    I13564,I13464,I13462,I24439,I24440,g23266,g13580,g10653,g11584,g16741,
    g13765,I14789,I14788,g19981,g13084,g12093,g14636,g12029,g12042,g11990,
    g11892,I17462,I17460,g17755,g14730,g14695,g16875,g14014,g16604,g12796,
    g27882,g14664,g13513,g13079,g13476,I22871,g12150,g13676,I22754,g24383,
    g28109,g12999,I22872,I22873,I14291,I14289,g11936,I15334,g12192,g10609,
    g22940,I12097,I12096,g25425,g20081,g12522,I22966,I22967,g17744,I17447,
    g13336,I17446,g17399,g12492,g15741,g34422,g9629,I13750,g12824,I12850,
    I12848,g11396,g8847,g11674,g8803,g15735,g14674,g11117,g7228,g10598,g29540,
    g22833,g21360,g12739,g12662,g13628,g14573,g14548,I15123,I15121,g12651,
    g10281,g17846,g14946,g17686,g17650,g16854,I29262,I29263,g10899,g11639,
    I13383,I13384,g7150,g10515,I25907,g26256,I20204,g26752,g25189,g11514,
    g16660,I26439,I26438,I29314,g14271,I23962,I12730,I12728,I12241,I12242,
    I29269,g12050,g14771,g12129,I12877,I12878,g11442,I13183,I13182,g12443,
    g17514,g12483,I15364,I15365,I14247,I15041,I13851,I13850,g24631,g23956,
    g12558,g12453,I32440,I32441,g12008,g16278,g8105,I23951,g13603,I23949,
    g26255,g24779,g12152,g16694,g17788,I29279,g12081,I29277,g15721,I29278,
    I14766,I14764,I15130,I15128,I15193,I29286,g12085,I29284,g12405,g11697,
    I14258,I14259,g13130,g11571,g19611,g13971,I12261,g12744,g12581,I18627,
    g14712,I18625,g26269,g26248,g17773,g17740,g14739,g16815,g13727,g15734,
    g20979,g23659,I13731,I13729,g31978,I22824,I22822,I15253,I18681,I18680,
    g13600,g11039,I22931,I22929,I20166,I20167,I15175,I15174,g34469,I32756,
    I14370,I14368,g26782,g25203,g11251,g11483,I15262,g22755,I12271,I12269,
    g13264,g11869,g24933,g19466,g7675,g13516,g11533,g11490,g11444,g11412,g9649,
    g14522,I31974,I31972,g12785,I15308,g13834,g13996,g22709,g22687,g9177,
    g11881,I29270,I29271,I18626,g12432,I22893,I22894,g23692,g20995,I26071,
    I26072,g11320,g24567,g22668,g19886,I15122,I14957,I14955,g22875,g13797,
    g11292,I14331,I14205,g9700,g12449,I14290,I22892,I14427,g14829,g12137,
    I31983,g14434,g11945,g9586,I12876,g10946,g12173,I13335,I13336,I11824,
    g14344,g11885,g22753,g22711,I17496,I17494,g14682,g12149,I14480,g12148,
    g13109,g16772,g13799,g24787,g23079,g13108,I22799,g11492,g12971,I12545,
    I12544,I13184,I14956,g27833,g14640,g17220,g9835,g17246,g12412,I26049,
    g13500,g12767,g22754,g33083,g12695,g13851,g13823,I22866,I22864,g21345,
    g9372,I20461,I20460,I12546,g24662,I24461,g14437,g15751,g13852,g12593,
    g12772,I26440,I22923,g21284,I22921,g29660,g14146,g14123,g16275,g13480,
    I14211,g12112,I17923,g13378,I14497,g14320,I24363,g13040,g12002,g8864,
    g27903,g12333,I12287,g14898,I32204,I32202,I23950,g24380,I23601,I23602,
    g14521,I25221,I17885,I17883,I13454,g22902,I16780,g12332,I16778,g9567,
    g24932,g15720,g14497,I14855,I14853,g29335,g25540,g28131,g13634,g24793,
    I12372,I24384,I24385,g13709,I18682,g17290,I29253,g12017,I15213,I15212,
    I12842,I14714,I14712,g22661,I13730,g27775,g13573,g13554,g13058,I14257,
    I15051,I14816,g22715,I23120,g14871,g14752,g12232,g16316,I22930,g12223,
    g17572,I14369,I22965,g12288,I32433,g24369,I23586,I23587,g10312,g21359,
    g10649,I13852,I12270,I14733,g17668,g17634,g17597,g14569,g21344,g16476,
    g12622,g10754,g11763,I12219,I12217,g25200,g23642,g12806,g11020,g12080,
    g13928,g11238,I12218,I20188,I20189,g29556,g24925,g20092,g17520,g12342,
    I22937,g12226,I22936,I26395,g14227,I26393,I14923,g12145,I15105,g13670,
    I23978,g21354,g10671,I16779,I12470,I12468,g9092,g10884,I12277,I13499,
    I13497,I17884,g12711,I12075,I12074,I26050,I26051,g24802,I23970,I23971,
    g15726,I13498,g23124,g26235,g24766,I14885,I14854,g12225,I15288,I15289,
    I29303,I29302,g14120,I22922,g14677,I25845,g26212,I15003,I15002,g13779,
    I22685,I26461,I23987,I23985,I22846,I12401,g27738,g16757,I20486,g13945,
    g16299,g8163,g17315,I23969,g14547,g12571,g13672,g16663,g14655,g23281,
    g22839,g23324,g20181,I20187,g21272,I13043,g17816,g17779,g11961,g12079,
    g13897,g11217,I24383,g14347,g12078,I26070,I11879,I11877,g12609,g13911,
    g13886,g11675,I11878,g12159,g12125,I21978,I21976,g24988,I15149,I15147,
    I23986,g24776,g26208,g16925,g14054,g16657,I15148,g27854,I26367,I26366,
    I26394,I15004,g13097,g13104,I15176,g14520,I14187,I25220,g16749,g13907,
    g33669,g10583,g7442,I13079,I13077,I32432,g14089,g22688,g16813,g13958,
    g16745,g13927,g17706,I13078,g14088,g17689,I18589,g14679,I18587,I18588,
    I20467,g16728,I14169,I14884,I17380,I17381,g12289,g12646,g14625,g14987,
    g17670,g13896,I23917,g23975,g25048,g26714,g11959,g11172,I22684,I12729,
    g13050,g20068,g14211,I14531,I14530,g13742,I14765,I12098,I12345,I14186,
    g14228,g12195,g17596,g12540,g17243,g14212,g12016,g21377,g14549,I18485,
    g14611,g15780,I17475,I17474,g14590,g12121,g12437,g25237,g22838,g17734,
    g13939,g9442,g25186,g26685,I15129,I26095,g11002,g12188,g12124,g11245,
    I14351,I14352,g21403,g17225,g12294,I18580,I18581,I11864,I14228,g17468,
    I21993,I21992,g14575,g14706,g17736,g14696,g17679,I14510,I14508,g15743,
    I13382,g22666,g13499,g11382,I13065,g11473,g13498,g12577,g12462,I15080,
    I15078,g17363,g14194,g21190,g17420,g12505,I23600,I14275,g12822,g12667,
    I15342,I24438,g14411,g15710,g9715,g10916,I12240,g12491,g12819,g12194,
    g13529,g11544,g11446,I14517,g12588,I26094,g12524,g20854,g13528,g13764,
    I12469,g12196,g9775,g9663,g12119,I22711,I22710,g15725,g15713,g12118,g15728,
    g13517,g16723,g13730,g22651,g11200,I24415,I24414,I15043,g13043,I17379,
    g13069,g13712,g15717,g13092,I13401,g11955,g11621,g19962,g10618,I14350,
    g25216,g34220,I18486,I18487,g14279,g12111,g9246,I12278,I12279,g15723,
    g10775,g13967,I14790,I12849,g22638,g14663,g8889,g10601,g13918,g14601,
    I18538,I12841,I15079,I12263,I14498,I14499,I15106,I15107,g20201,I20468,
    I20469,g22405,g13086,g17578,g7167,g10537,g12185,g17757,g14740,g17716,
    g14638,g11977,g34227,I32203,g25172,g23560,g16687,g11858,I17405,g25019,
    g15742,g9203,I13518,g29497,g12083,g14556,g14382,I29261,g12046,g19965,
    g24808,g17571,g7304,g9509,g15709,I25243,g13518,I14509,I13566,I22793,g10928,
    g13240,g13115,g8227,g12115,I13139,g13544,g24570,I15042,I15255,g11189,
    I14248,I14249,g23210,g16696,g13871,g13882,g10578,g11938,g12371,I32518,
    g13908,g17364,g12207,I12262,I14213,g15736,g17635,I17448,I22945,g14517,
    g25175,g17708,g17640,g14598,I32439,g22713,I14428,I14429,g11155,g13083,
    g13822,I15167,I22823,g14600,g14781,g24576,g21417,I14170,I14171,g12114,
    g13118,g22850,g22650,I20462,I21977,I22900,I22901,I15053,I15254,I25846,
    I25847,g14422,g16770,g22757,g20055,g20107,g14542,g21283,I22865,g10614,
    g12049,g17775,I17925,g11914,g17872,g14602,g7184,g10561,g11924,g7209,g13910,
    g19632,I14212,I18531,I17924,I29255,g17820,I29285,g15752,I13463,g17396,
    g14272,g14750,I14713,I17461,I12076,g19916,g23105,g13139,g21253,g17482,
    I22938,g15729,g13098,g26666,g25144,g21331,I15052,I14925,I17495,I26368,
    g24951,g13798,g11973,g23726,g21140,g25160,g14574,g14452,I17476,g17647,
    I14610,I14611,g20163,g15782,I29254,I15214,g12045,g17513,g13241,g23602,
    I22712,g10929,g23756,g17723,g17495,g13515,g12628,I23918,I23919,g23678,
    I14276,I14277,g13883,g14803,g10737,g12147,I14924,g22837,g12151,I20223,
    g27377,I21994,g16313,g12227,I31973,I29304,g14678,I18579,g13970,g12044,
    g17765,g20172,g23357,g12120,g23711,g10961,g16424,g11216,g12189,g12146,
    g21206,g24751,g23052,I24416,I14532,g19442,g25381,g17598,g8131,g11173,
    g12190,g29503,g11231,g11907,g11134,g19887,g10603,g15798,g11903,g11862,
    g8347,g22643,I13066,I13067,g17792,g12479,g13462,g10611,g11107,g24943,
    g11248,g15788,g12287,g17669,g17309,g13551,g17705,I12253,g15829,g13831,
    g19913,g10336,g12486,g12252,g12166,g15718,g10488,g16220,g23955,g12123,
    g23918,g13661,g12821,g10555,g16581,g22190,g23686,g19778,g16232,g23051,
    g19793,g8086,g11363,g16231,g13622,g23883,g16201,g16210,g12204,g16242,
    g16209,g12364,g19853,g14792,g15724,g12970,g10510,g23871,g11309,g12314,
    g19873,g12435,g10179,g23024,g23763,g11276,g16219,g14751,g31294,g10205,
    g23835,g16488;

  FD1 DFF_0(CK,g5057,g33046);
  FD1 DFF_1(CK,g2771,g34441);
  FD1 DFF_2(CK,g1882,g33982);
  FD1 DFF_3(CK,g6462,g25751);
  FD1 DFF_4(CK,g2299,g34007);
  FD1 DFF_5(CK,g4040,g24276);
  FD1 DFF_6(CK,g2547,g30381);
  FD1 DFF_7(CK,g559,g640);
  FD1 DFF_8(CK,g3017,g31877);
  FD1 DFF_9(CK,g3243,g30405);
  FD1 DFF_10(CK,g452,g25604);
  FD1 DFF_11(CK,g464,g25607);
  FD1 DFF_12(CK,g3542,g30416);
  FD1 DFF_13(CK,g5232,g30466);
  FD1 DFF_14(CK,g5813,g25736);
  FD1 DFF_15(CK,g2907,g34617);
  FD1 DFF_16(CK,g1744,g33974);
  FD1 DFF_17(CK,g5909,g30505);
  FD1 DFF_18(CK,g1802,g33554);
  FD1 DFF_19(CK,g3554,g30432);
  FD1 DFF_20(CK,g6219,g33064);
  FD1 DFF_21(CK,g807,g34881);
  FD1 DFF_22(CK,g6031,g6027);
  FD1 DFF_23(CK,g847,g24216);
  FD1 DFF_24(CK,g976,g24232);
  FD1 DFF_25(CK,g4172,g34733);
  FD1 DFF_26(CK,g4372,g34882);
  FD1 DFF_27(CK,g3512,g33026);
  FD1 DFF_28(CK,g749,g31867);
  FD1 DFF_29(CK,g3490,g25668);
  FD1 DFF_30(CK,g6005,g24344);
  FD1 DFF_31(CK,g4235,g4232);
  FD1 DFF_32(CK,g1600,g33966);
  FD1 DFF_33(CK,g1714,g33550);
  FD1 DFF_34(CK,g3649,g3625);
  FD1 DFF_35(CK,g3155,g30393);
  FD1 DFF_36(CK,g3355,g31880);
  FD1 DFF_37(CK,g2236,g29248);
  FD1 DFF_38(CK,g4555,g4571);
  FD1 DFF_39(CK,g3698,g24274);
  FD1 DFF_40(CK,g6073,g31920);
  FD1 DFF_41(CK,g1736,g33973);
  FD1 DFF_42(CK,g1968,g30360);
  FD1 DFF_43(CK,g4621,g34460);
  FD1 DFF_44(CK,g5607,g30494);
  FD1 DFF_45(CK,g2657,g30384);
  FD1 DFF_46(CK,g5659,g24340);
  FD1 DFF_47(CK,g490,g29223);
  FD1 DFF_48(CK,g311,g26881);
  FD1 DFF_49(CK,g6069,g31925);
  FD1 DFF_50(CK,g772,g34252);
  FD1 DFF_51(CK,g5587,g30489);
  FD1 DFF_52(CK,g6177,g29301);
  FD1 DFF_53(CK,g6377,g6373);
  FD1 DFF_54(CK,g3167,g33022);
  FD1 DFF_55(CK,g5615,g30496);
  FD1 DFF_56(CK,g4567,g33043);
  FD1 DFF_57(CK,g3057,g28062);
  FD1 DFF_58(CK,g3457,g29263);
  FD1 DFF_59(CK,g6287,g30533);
  FD1 DFF_60(CK,g1500,g24256);
  FD1 DFF_61(CK,g2563,g34015);
  FD1 DFF_62(CK,g4776,g34031);
  FD1 DFF_63(CK,g4593,g34452);
  FD1 DFF_64(CK,g6199,g34646);
  FD1 DFF_65(CK,g2295,g34001);
  FD1 DFF_66(CK,g1384,g25633);
  FD1 DFF_67(CK,g1339,g24259);
  FD1 DFF_68(CK,g5180,g33049);
  FD1 DFF_69(CK,g2844,g34609);
  FD1 DFF_70(CK,g1024,g31869);
  FD1 DFF_71(CK,g5591,g30490);
  FD1 DFF_72(CK,g3598,g30427);
  FD1 DFF_73(CK,g4264,g21894);
  FD1 DFF_74(CK,g767,g33965);
  FD1 DFF_75(CK,g5853,g34645);
  FD1 DFF_76(CK,g3321,g3317);
  FD1 DFF_77(CK,g2089,g33571);
  FD1 DFF_78(CK,g4933,g34267);
  FD1 DFF_79(CK,g4521,g26971);
  FD1 DFF_80(CK,g5507,g34644);
  FD1 DFF_81(CK,g3625,g3618);
  FD1 DFF_82(CK,g6291,g30534);
  FD1 DFF_83(CK,g294,g33535);
  FD1 DFF_84(CK,g5559,g30498);
  FD1 DFF_85(CK,g5794,g25728);
  FD1 DFF_86(CK,g6144,g25743);
  FD1 DFF_87(CK,g3813,g25684);
  FD1 DFF_88(CK,g562,g25613);
  FD1 DFF_89(CK,g608,g34438);
  FD1 DFF_90(CK,g1205,g24244);
  FD1 DFF_91(CK,g3909,g30439);
  FD1 DFF_92(CK,g6259,g30541);
  FD1 DFF_93(CK,g5905,g30519);
  FD1 DFF_94(CK,g921,g25621);
  FD1 DFF_95(CK,g2955,g34807);
  FD1 DFF_96(CK,g203,g25599);
  FD1 DFF_97(CK,g6088,g31924);
  FD1 DFF_98(CK,g1099,g24235);
  FD1 DFF_99(CK,g4878,g34036);
  FD1 DFF_100(CK,g5204,g30476);
  FD1 DFF_101(CK,g5630,g5623);
  FD1 DFF_102(CK,g3606,g30429);
  FD1 DFF_103(CK,g1926,g32997);
  FD1 DFF_104(CK,g6215,g33063);
  FD1 DFF_105(CK,g3586,g30424);
  FD1 DFF_106(CK,g291,g32977);
  FD1 DFF_107(CK,g4674,g34026);
  FD1 DFF_108(CK,g3570,g30420);
  FD1 DFF_109(CK,g640,g637);
  FD1 DFF_110(CK,g5969,g6012);
  FD1 DFF_111(CK,g1862,g33560);
  FD1 DFF_112(CK,g676,g29226);
  FD1 DFF_113(CK,g843,g25619);
  FD1 DFF_114(CK,g4132,g28076);
  FD1 DFF_115(CK,g4332,g34455);
  FD1 DFF_116(CK,g4153,g30457);
  FD1 DFF_117(CK,g5666,g5637);
  FD1 DFF_118(CK,g6336,g33625);
  FD1 DFF_119(CK,g622,g34790);
  FD1 DFF_120(CK,g3506,g30414);
  FD1 DFF_121(CK,g4558,g26966);
  FD1 DFF_122(CK,g6065,g31923);
  FD1 DFF_123(CK,g6322,g6315);
  FD1 DFF_124(CK,g3111,g25656);
  FD1 DFF_125(CK,g117,g30390);
  FD1 DFF_126(CK,g2837,g26935);
  FD1 DFF_127(CK,g939,g34727);
  FD1 DFF_128(CK,g278,g25594);
  FD1 DFF_129(CK,g4492,g26963);
  FD1 DFF_130(CK,g4864,g34034);
  FD1 DFF_131(CK,g1036,g33541);
  FD1 DFF_132(CK,g128,g28093);
  FD1 DFF_133(CK,g1178,g24236);
  FD1 DFF_134(CK,g3239,g30404);
  FD1 DFF_135(CK,g718,g28051);
  FD1 DFF_136(CK,g6195,g29303);
  FD1 DFF_137(CK,g1135,g26917);
  FD1 DFF_138(CK,g6137,g25741);
  FD1 DFF_139(CK,g6395,g33624);
  FD1 DFF_140(CK,g3380,g31882);
  FD1 DFF_141(CK,g5343,g24337);
  FD1 DFF_142(CK,g554,g34911);
  FD1 DFF_143(CK,g496,g33963);
  FD1 DFF_144(CK,g3853,g34627);
  FD1 DFF_145(CK,g5134,g29282);
  FD1 DFF_146(CK,g1422,g1418);
  FD1 DFF_147(CK,g3794,g25676);
  FD1 DFF_148(CK,g2485,g33013);
  FD1 DFF_149(CK,g925,g32981);
  FD1 DFF_150(CK,g48,g34993);
  FD1 DFF_151(CK,g5555,g30483);
  FD1 DFF_152(CK,g878,g875);
  FD1 DFF_153(CK,g1798,g32994);
  FD1 DFF_154(CK,g4076,g28070);
  FD1 DFF_155(CK,g2941,g34806);
  FD1 DFF_156(CK,g3905,g30453);
  FD1 DFF_157(CK,g763,g33539);
  FD1 DFF_158(CK,g6255,g30526);
  FD1 DFF_159(CK,g4375,g26951);
  FD1 DFF_160(CK,g4871,g34035);
  FD1 DFF_161(CK,g4722,g34636);
  FD1 DFF_162(CK,g590,g32978);
  FD1 DFF_163(CK,g6692,g6668);
  FD1 DFF_164(CK,g1632,g30348);
  FD1 DFF_165(CK,g5313,g24336);
  FD1 DFF_166(CK,g3100,g3092);
  FD1 DFF_167(CK,g1495,g24250);
  FD1 DFF_168(CK,g6497,g6490);
  FD1 DFF_169(CK,g1437,g29236);
  FD1 DFF_170(CK,g6154,g29298);
  FD1 DFF_171(CK,g1579,g1576);
  FD1 DFF_172(CK,g5567,g30499);
  FD1 DFF_173(CK,g1752,g33976);
  FD1 DFF_174(CK,g1917,g32996);
  FD1 DFF_175(CK,g744,g30335);
  FD1 DFF_176(CK,g3040,g31878);
  FD1 DFF_177(CK,g4737,g34637);
  FD1 DFF_178(CK,g4809,g25693);
  FD1 DFF_179(CK,g6267,g30528);
  FD1 DFF_180(CK,g3440,g25661);
  FD1 DFF_181(CK,g3969,g4012);
  FD1 DFF_182(CK,g1442,g24251);
  FD1 DFF_183(CK,g5965,g30521);
  FD1 DFF_184(CK,g4477,g26960);
  FD1 DFF_185(CK,g1233,g24239);
  FD1 DFF_186(CK,g4643,g34259);
  FD1 DFF_187(CK,g5264,g30474);
  FD1 DFF_188(CK,g6329,g6351);
  FD1 DFF_189(CK,g2610,g33016);
  FD1 DFF_190(CK,g5160,g34643);
  FD1 DFF_191(CK,g5360,g31905);
  FD1 DFF_192(CK,g5933,g30510);
  FD1 DFF_193(CK,g1454,g29239);
  FD1 DFF_194(CK,g753,g26897);
  FD1 DFF_195(CK,g1296,g34729);
  FD1 DFF_196(CK,g3151,g34625);
  FD1 DFF_197(CK,g2980,g34800);
  FD1 DFF_198(CK,g6727,g24353);
  FD1 DFF_199(CK,g3530,g33029);
  FD1 DFF_200(CK,g4742,g21903);
  FD1 DFF_201(CK,g4104,g33615);
  FD1 DFF_202(CK,g1532,g24253);
  FD1 DFF_203(CK,g4304,g24281);
  FD1 DFF_204(CK,g2177,g33997);
  FD1 DFF_205(CK,g3010,g25651);
  FD1 DFF_206(CK,g52,g34997);
  FD1 DFF_207(CK,g4754,g34263);
  FD1 DFF_208(CK,g1189,g24237);
  FD1 DFF_209(CK,g2287,g33584);
  FD1 DFF_210(CK,g4273,g24280);
  FD1 DFF_211(CK,g1389,g26920);
  FD1 DFF_212(CK,g1706,g33548);
  FD1 DFF_213(CK,g5835,g29296);
  FD1 DFF_214(CK,g1171,g30338);
  FD1 DFF_215(CK,g4269,g21895);
  FD1 DFF_216(CK,g2399,g33588);
  FD1 DFF_217(CK,g3372,g31886);
  FD1 DFF_218(CK,g4983,g34041);
  FD1 DFF_219(CK,g5611,g30495);
  FD1 DFF_220(CK,g3618,g3661);
  FD1 DFF_221(CK,g4572,g29279);
  FD1 DFF_222(CK,g3143,g25655);
  FD1 DFF_223(CK,g2898,g34795);
  FD1 DFF_224(CK,g3343,g24269);
  FD1 DFF_225(CK,g3235,g30403);
  FD1 DFF_226(CK,g4543,g33042);
  FD1 DFF_227(CK,g3566,g30419);
  FD1 DFF_228(CK,g4534,g34023);
  FD1 DFF_229(CK,g4961,g28090);
  FD1 DFF_230(CK,g6398,g31926);
  FD1 DFF_231(CK,g4927,g34642);
  FD1 DFF_232(CK,g2259,g30370);
  FD1 DFF_233(CK,g2819,g34448);
  FD1 DFF_234(CK,g4414,g26946);
  FD1 DFF_235(CK,g5802,g5794);
  FD1 DFF_236(CK,g2852,g34610);
  FD1 DFF_237(CK,g417,g24209);
  FD1 DFF_238(CK,g681,g28047);
  FD1 DFF_239(CK,g437,g24206);
  FD1 DFF_240(CK,g351,g26891);
  FD1 DFF_241(CK,g5901,g30504);
  FD1 DFF_242(CK,g2886,g34798);
  FD1 DFF_243(CK,g3494,g25669);
  FD1 DFF_244(CK,g5511,g30480);
  FD1 DFF_245(CK,g3518,g33027);
  FD1 DFF_246(CK,g1604,g33972);
  FD1 DFF_247(CK,g4135,g28077);
  FD1 DFF_248(CK,g5092,g25697);
  FD1 DFF_249(CK,g4831,g28099);
  FD1 DFF_250(CK,g4382,g26947);
  FD1 DFF_251(CK,g6386,g24350);
  FD1 DFF_252(CK,g479,g24210);
  FD1 DFF_253(CK,g3965,g30455);
  FD1 DFF_254(CK,g4749,g28084);
  FD1 DFF_255(CK,g2008,g33993);
  FD1 DFF_256(CK,g736,g802);
  FD1 DFF_257(CK,g3933,g30444);
  FD1 DFF_258(CK,g222,g33537);
  FD1 DFF_259(CK,g3050,g25650);
  FD1 DFF_260(CK,g5736,g31915);
  FD1 DFF_261(CK,g1052,g25625);
  FD1 DFF_262(CK,g58,g30328);
  FD1 DFF_263(CK,g5623,g5666);
  FD1 DFF_264(CK,g2122,g30366);
  FD1 DFF_265(CK,g2465,g33593);
  FD1 DFF_266(CK,g6483,g25755);
  FD1 DFF_267(CK,g5889,g30502);
  FD1 DFF_268(CK,g4495,g33036);
  FD1 DFF_269(CK,g365,g25595);
  FD1 DFF_270(CK,g4653,g34462);
  FD1 DFF_271(CK,g3179,g33024);
  FD1 DFF_272(CK,g1728,g33552);
  FD1 DFF_273(CK,g2433,g34014);
  FD1 DFF_274(CK,g3835,g29273);
  FD1 DFF_275(CK,g6187,g25748);
  FD1 DFF_276(CK,g4917,g34638);
  FD1 DFF_277(CK,g1070,g30341);
  FD1 DFF_278(CK,g822,g26899);
  FD1 DFF_279(CK,g6027,g6023);
  FD1 DFF_280(CK,g914,g30336);
  FD1 DFF_281(CK,g5339,g5335);
  FD1 DFF_282(CK,g4164,g26940);
  FD1 DFF_283(CK,g969,g25622);
  FD1 DFF_284(CK,g2807,g34447);
  FD1 DFF_285(CK,g5424,g25709);
  FD1 DFF_286(CK,g4054,g33613);
  FD1 DFF_287(CK,g6191,g25749);
  FD1 DFF_288(CK,g5077,g25704);
  FD1 DFF_289(CK,g5523,g33053);
  FD1 DFF_290(CK,g3680,g3676);
  FD1 DFF_291(CK,g6637,g30555);
  FD1 DFF_292(CK,g174,g25601);
  FD1 DFF_293(CK,g1682,g33971);
  FD1 DFF_294(CK,g355,g26892);
  FD1 DFF_295(CK,g1087,g1083);
  FD1 DFF_296(CK,g1105,g26915);
  FD1 DFF_297(CK,g2342,g33008);
  FD1 DFF_298(CK,g6307,g30538);
  FD1 DFF_299(CK,g3802,g3794);
  FD1 DFF_300(CK,g6159,g25750);
  FD1 DFF_301(CK,g2255,g30369);
  FD1 DFF_302(CK,g2815,g34446);
  FD1 DFF_303(CK,g911,g29230);
  FD1 DFF_304(CK,g43,g34789);
  FD1 DFF_305(CK,g4012,g3983);
  FD1 DFF_306(CK,g1748,g33975);
  FD1 DFF_307(CK,g5551,g30497);
  FD1 DFF_308(CK,g5742,g31917);
  FD1 DFF_309(CK,g3558,g30418);
  FD1 DFF_310(CK,g5499,g25721);
  FD1 DFF_311(CK,g2960,g34622);
  FD1 DFF_312(CK,g3901,g30438);
  FD1 DFF_313(CK,g4888,g34266);
  FD1 DFF_314(CK,g6251,g30540);
  FD1 DFF_315(CK,g6315,g6358);
  FD1 DFF_316(CK,g1373,g32986);
  FD1 DFF_317(CK,g3092,g25648);
  FD1 DFF_318(CK,g157,g33960);
  FD1 DFF_319(CK,g2783,g34442);
  FD1 DFF_320(CK,g4281,g4277);
  FD1 DFF_321(CK,g3574,g30421);
  FD1 DFF_322(CK,g2112,g33573);
  FD1 DFF_323(CK,g1283,g34730);
  FD1 DFF_324(CK,g433,g24205);
  FD1 DFF_325(CK,g4297,g4294);
  FD1 DFF_326(CK,g5983,g6005);
  FD1 DFF_327(CK,g1459,g1399);
  FD1 DFF_328(CK,g758,g32979);
  FD1 DFF_329(CK,g5712,g25731);
  FD1 DFF_330(CK,g4138,g28078);
  FD1 DFF_331(CK,g4639,g34025);
  FD1 DFF_332(CK,g6537,g25763);
  FD1 DFF_333(CK,g5543,g30481);
  FD1 DFF_334(CK,g1582,g1500);
  FD1 DFF_335(CK,g3736,g31890);
  FD1 DFF_336(CK,g5961,g30517);
  FD1 DFF_337(CK,g6243,g30539);
  FD1 DFF_338(CK,g632,g34880);
  FD1 DFF_339(CK,g1227,g24242);
  FD1 DFF_340(CK,g3889,g30436);
  FD1 DFF_341(CK,g3476,g29265);
  FD1 DFF_342(CK,g1664,g32990);
  FD1 DFF_343(CK,g1246,g24245);
  FD1 DFF_344(CK,g6128,g25739);
  FD1 DFF_345(CK,g6629,g30553);
  FD1 DFF_346(CK,g246,g26907);
  FD1 DFF_347(CK,g4049,g24278);
  FD1 DFF_348(CK,g4449,g26955);
  FD1 DFF_349(CK,g2932,g24282);
  FD1 DFF_350(CK,g4575,g29276);
  FD1 DFF_351(CK,g4098,g31894);
  FD1 DFF_352(CK,g4498,g33037);
  FD1 DFF_353(CK,g528,g26894);
  FD1 DFF_354(CK,g5436,g25711);
  FD1 DFF_355(CK,g16,g34593);
  FD1 DFF_356(CK,g3139,g25654);
  FD1 DFF_357(CK,g102,g33962);
  FD1 DFF_358(CK,g4584,g34451);
  FD1 DFF_359(CK,g142,g34250);
  FD1 DFF_360(CK,g5335,g5331);
  FD1 DFF_361(CK,g5831,g29295);
  FD1 DFF_362(CK,g239,g26905);
  FD1 DFF_363(CK,g1216,g25629);
  FD1 DFF_364(CK,g2848,g34792);
  FD1 DFF_365(CK,g5805,g5798);
  FD1 DFF_366(CK,g5022,g25703);
  FD1 DFF_367(CK,g4019,g4000);
  FD1 DFF_368(CK,g1030,g32983);
  FD1 DFF_369(CK,g3672,g3668);
  FD1 DFF_370(CK,g3231,g30402);
  FD1 DFF_371(CK,g6490,g25757);
  FD1 DFF_372(CK,g1430,g1426);
  FD1 DFF_373(CK,g4452,g4446);
  FD1 DFF_374(CK,g2241,g33999);
  FD1 DFF_375(CK,g1564,g24262);
  FD1 DFF_376(CK,g5798,g25729);
  FD1 DFF_377(CK,g6148,g6140);
  FD1 DFF_378(CK,g6649,g30558);
  FD1 DFF_379(CK,g110,g34848);
  FD1 DFF_380(CK,g884,g881);
  FD1 DFF_381(CK,g3742,g31892);
  FD1 DFF_382(CK,g225,g26901);
  FD1 DFF_383(CK,g4486,g26961);
  FD1 DFF_384(CK,g4504,g33039);
  FD1 DFF_385(CK,g5873,g33059);
  FD1 DFF_386(CK,g5037,g31899);
  FD1 DFF_387(CK,g2319,g33007);
  FD1 DFF_388(CK,g5495,g25720);
  FD1 DFF_389(CK,g4185,g21891);
  FD1 DFF_390(CK,g5208,g30462);
  FD1 DFF_391(CK,g2152,g18422);
  FD1 DFF_392(CK,g5579,g30487);
  FD1 DFF_393(CK,g5869,g33058);
  FD1 DFF_394(CK,g5719,g31916);
  FD1 DFF_395(CK,g1589,g24261);
  FD1 DFF_396(CK,g5752,g25730);
  FD1 DFF_397(CK,g6279,g30531);
  FD1 DFF_398(CK,g5917,g30506);
  FD1 DFF_399(CK,g2975,g34804);
  FD1 DFF_400(CK,g6167,g25747);
  FD1 DFF_401(CK,g3983,g4005);
  FD1 DFF_402(CK,g2599,g33601);
  FD1 DFF_403(CK,g1448,g26922);
  FD1 DFF_404(CK,g881,g878);
  FD1 DFF_405(CK,g3712,g25679);
  FD1 DFF_406(CK,g2370,g29250);
  FD1 DFF_407(CK,g5164,g30459);
  FD1 DFF_408(CK,g1333,g1582);
  FD1 DFF_409(CK,g153,g33534);
  FD1 DFF_410(CK,g6549,g30543);
  FD1 DFF_411(CK,g4087,g29275);
  FD1 DFF_412(CK,g4801,g34030);
  FD1 DFF_413(CK,g2984,g34980);
  FD1 DFF_414(CK,g3961,g30451);
  FD1 DFF_415(CK,g5770,g25723);
  FD1 DFF_416(CK,g962,g25627);
  FD1 DFF_417(CK,g101,g34787);
  FD1 DFF_418(CK,g4226,g4222);
  FD1 DFF_419(CK,g6625,g30552);
  FD1 DFF_420(CK,g51,g34996);
  FD1 DFF_421(CK,g1018,g30337);
  FD1 DFF_422(CK,g1418,g24254);
  FD1 DFF_423(CK,g4045,g24277);
  FD1 DFF_424(CK,g1467,g29237);
  FD1 DFF_425(CK,g2461,g30378);
  FD1 DFF_426(CK,g5706,g31912);
  FD1 DFF_427(CK,g457,g25603);
  FD1 DFF_428(CK,g2756,g33019);
  FD1 DFF_429(CK,g5990,g33623);
  FD1 DFF_430(CK,g471,g25608);
  FD1 DFF_431(CK,g1256,g29235);
  FD1 DFF_432(CK,g5029,g31902);
  FD1 DFF_433(CK,g6519,g29306);
  FD1 DFF_434(CK,g4169,g28080);
  FD1 DFF_435(CK,g1816,g33978);
  FD1 DFF_436(CK,g4369,g26970);
  FD1 DFF_437(CK,g3436,g25660);
  FD1 DFF_438(CK,g5787,g25726);
  FD1 DFF_439(CK,g4578,g29278);
  FD1 DFF_440(CK,g4459,g34253);
  FD1 DFF_441(CK,g3831,g29272);
  FD1 DFF_442(CK,g2514,g33595);
  FD1 DFF_443(CK,g3288,g33610);
  FD1 DFF_444(CK,g2403,g33589);
  FD1 DFF_445(CK,g2145,g34605);
  FD1 DFF_446(CK,g1700,g30350);
  FD1 DFF_447(CK,g513,g25611);
  FD1 DFF_448(CK,g2841,g26936);
  FD1 DFF_449(CK,g5297,g33619);
  FD1 DFF_450(CK,g3805,g3798);
  FD1 DFF_451(CK,g2763,g34022);
  FD1 DFF_452(CK,g4793,g34033);
  FD1 DFF_453(CK,g952,g34726);
  FD1 DFF_454(CK,g1263,g31870);
  FD1 DFF_455(CK,g1950,g33985);
  FD1 DFF_456(CK,g5138,g29283);
  FD1 DFF_457(CK,g2307,g34003);
  FD1 DFF_458(CK,g5109,g5101);
  FD1 DFF_459(CK,g5791,g25727);
  FD1 DFF_460(CK,g3798,g25677);
  FD1 DFF_461(CK,g4664,g34463);
  FD1 DFF_462(CK,g2223,g33006);
  FD1 DFF_463(CK,g5808,g29292);
  FD1 DFF_464(CK,g6645,g30557);
  FD1 DFF_465(CK,g2016,g33989);
  FD1 DFF_466(CK,g5759,g28098);
  FD1 DFF_467(CK,g3873,g33033);
  FD1 DFF_468(CK,g3632,g3654);
  FD1 DFF_469(CK,g2315,g34005);
  FD1 DFF_470(CK,g2811,g26932);
  FD1 DFF_471(CK,g5957,g30516);
  FD1 DFF_472(CK,g2047,g33575);
  FD1 DFF_473(CK,g3869,g33032);
  FD1 DFF_474(CK,g6358,g6329);
  FD1 DFF_475(CK,g3719,g31891);
  FD1 DFF_476(CK,g5575,g30486);
  FD1 DFF_477(CK,g46,g34991);
  FD1 DFF_478(CK,g3752,g25678);
  FD1 DFF_479(CK,g3917,g30440);
  FD1 DFF_480(CK,g4188,g4191);
  FD1 DFF_481(CK,g1585,g1570);
  FD1 DFF_482(CK,g4388,g26949);
  FD1 DFF_483(CK,g6275,g30530);
  FD1 DFF_484(CK,g6311,g30542);
  FD1 DFF_485(CK,g4216,g4213);
  FD1 DFF_486(CK,g1041,g25624);
  FD1 DFF_487(CK,g2595,g30383);
  FD1 DFF_488(CK,g2537,g33597);
  FD1 DFF_489(CK,g136,g34598);
  FD1 DFF_490(CK,g4430,g26957);
  FD1 DFF_491(CK,g4564,g26967);
  FD1 DFF_492(CK,g3454,g3447);
  FD1 DFF_493(CK,g4826,g28102);
  FD1 DFF_494(CK,g6239,g30524);
  FD1 DFF_495(CK,g3770,g25671);
  FD1 DFF_496(CK,g232,g26903);
  FD1 DFF_497(CK,g5268,g30475);
  FD1 DFF_498(CK,g6545,g34647);
  FD1 DFF_499(CK,g2417,g30377);
  FD1 DFF_500(CK,g1772,g33553);
  FD1 DFF_501(CK,g4741,g21902);
  FD1 DFF_502(CK,g5052,g31903);
  FD1 DFF_503(CK,g5452,g25715);
  FD1 DFF_504(CK,g1890,g33984);
  FD1 DFF_505(CK,g2629,g33602);
  FD1 DFF_506(CK,g572,g28045);
  FD1 DFF_507(CK,g2130,g34603);
  FD1 DFF_508(CK,g4108,g33035);
  FD1 DFF_509(CK,g4308,g4304);
  FD1 DFF_510(CK,g475,g24208);
  FD1 DFF_511(CK,g990,g1239);
  FD1 DFF_512(CK,g31,g34596);
  FD1 DFF_513(CK,g3412,g28064);
  FD1 DFF_514(CK,g45,g34990);
  FD1 DFF_515(CK,g799,g24213);
  FD1 DFF_516(CK,g3706,g31887);
  FD1 DFF_517(CK,g3990,g33614);
  FD1 DFF_518(CK,g5385,g31907);
  FD1 DFF_519(CK,g5881,g33060);
  FD1 DFF_520(CK,g1992,g30362);
  FD1 DFF_521(CK,g3029,g31875);
  FD1 DFF_522(CK,g3171,g33023);
  FD1 DFF_523(CK,g3787,g25674);
  FD1 DFF_524(CK,g812,g26898);
  FD1 DFF_525(CK,g832,g25618);
  FD1 DFF_526(CK,g5897,g30518);
  FD1 DFF_527(CK,g4165,g28079);
  FD1 DFF_528(CK,g4571,g6974);
  FD1 DFF_529(CK,g3281,g3303);
  FD1 DFF_530(CK,g4455,g26959);
  FD1 DFF_531(CK,g2902,g34801);
  FD1 DFF_532(CK,g333,g26884);
  FD1 DFF_533(CK,g168,g25600);
  FD1 DFF_534(CK,g2823,g26933);
  FD1 DFF_535(CK,g3684,g28066);
  FD1 DFF_536(CK,g3639,g33612);
  FD1 DFF_537(CK,g5331,g5327);
  FD1 DFF_538(CK,g3338,g24268);
  FD1 DFF_539(CK,g5406,g25716);
  FD1 DFF_540(CK,g3791,g25675);
  FD1 DFF_541(CK,g269,g26906);
  FD1 DFF_542(CK,g401,g24203);
  FD1 DFF_543(CK,g6040,g24346);
  FD1 DFF_544(CK,g441,g24207);
  FD1 DFF_545(CK,g5105,g25701);
  FD1 DFF_546(CK,g3808,g29269);
  FD1 DFF_547(CK,g9,g34592);
  FD1 DFF_548(CK,g3759,g28068);
  FD1 DFF_549(CK,g4467,g34255);
  FD1 DFF_550(CK,g3957,g30450);
  FD1 DFF_551(CK,g4093,g30456);
  FD1 DFF_552(CK,g1760,g32991);
  FD1 DFF_553(CK,g6151,g6144);
  FD1 DFF_554(CK,g6351,g24348);
  FD1 DFF_555(CK,g160,g34249);
  FD1 DFF_556(CK,g5445,g25713);
  FD1 DFF_557(CK,g5373,g31909);
  FD1 DFF_558(CK,g2279,g30371);
  FD1 DFF_559(CK,g3498,g29268);
  FD1 DFF_560(CK,g586,g29224);
  FD1 DFF_561(CK,g869,g859);
  FD1 DFF_562(CK,g2619,g33017);
  FD1 DFF_563(CK,g1183,g30339);
  FD1 DFF_564(CK,g1608,g33967);
  FD1 DFF_565(CK,g4197,g4194);
  FD1 DFF_566(CK,g5283,g5276);
  FD1 DFF_567(CK,g1779,g33559);
  FD1 DFF_568(CK,g2652,g29255);
  FD1 DFF_569(CK,g5459,g5452);
  FD1 DFF_570(CK,g2193,g30368);
  FD1 DFF_571(CK,g2393,g30375);
  FD1 DFF_572(CK,g5767,g25732);
  FD1 DFF_573(CK,g661,g28052);
  FD1 DFF_574(CK,g4950,g28089);
  FD1 DFF_575(CK,g5535,g33055);
  FD1 DFF_576(CK,g2834,g30392);
  FD1 DFF_577(CK,g1361,g30343);
  FD1 DFF_578(CK,g3419,g25657);
  FD1 DFF_579(CK,g6235,g30523);
  FD1 DFF_580(CK,g1146,g24233);
  FD1 DFF_581(CK,g2625,g33018);
  FD1 DFF_582(CK,g150,g32976);
  FD1 DFF_583(CK,g1696,g30349);
  FD1 DFF_584(CK,g6555,g33067);
  FD1 DFF_585(CK,g859,g26900);
  FD1 DFF_586(CK,g3385,g31883);
  FD1 DFF_587(CK,g3881,g33034);
  FD1 DFF_588(CK,g6621,g30551);
  FD1 DFF_589(CK,g3470,g25667);
  FD1 DFF_590(CK,g3897,g30452);
  FD1 DFF_591(CK,g518,g25612);
  FD1 DFF_592(CK,g3025,g31874);
  FD1 DFF_593(CK,g538,g34719);
  FD1 DFF_594(CK,g2606,g33607);
  FD1 DFF_595(CK,g1472,g26923);
  FD1 DFF_596(CK,g6113,g25746);
  FD1 DFF_597(CK,g542,g24211);
  FD1 DFF_598(CK,g5188,g33050);
  FD1 DFF_599(CK,g5689,g24341);
  FD1 DFF_600(CK,g1116,g1056);
  FD1 DFF_601(CK,g405,g24201);
  FD1 DFF_602(CK,g5216,g30463);
  FD1 DFF_603(CK,g6494,g6486);
  FD1 DFF_604(CK,g4669,g34464);
  FD1 DFF_605(CK,g5428,g25710);
  FD1 DFF_606(CK,g996,g24243);
  FD1 DFF_607(CK,g4531,g24335);
  FD1 DFF_608(CK,g2860,g34611);
  FD1 DFF_609(CK,g4743,g34262);
  FD1 DFF_610(CK,g6593,g30546);
  FD1 DFF_611(CK,g2710,g18527);
  FD1 DFF_612(CK,g215,g25591);
  FD1 DFF_613(CK,g4411,g4414);
  FD1 DFF_614(CK,g1413,g30347);
  FD1 DFF_615(CK,g4474,g10384);
  FD1 DFF_616(CK,g5308,g5283);
  FD1 DFF_617(CK,g6641,g30556);
  FD1 DFF_618(CK,g3045,g33020);
  FD1 DFF_619(CK,g6,g34589);
  FD1 DFF_620(CK,g1936,g33562);
  FD1 DFF_621(CK,g55,g35002);
  FD1 DFF_622(CK,g504,g25610);
  FD1 DFF_623(CK,g2587,g33015);
  FD1 DFF_624(CK,g4480,g31896);
  FD1 DFF_625(CK,g2311,g34004);
  FD1 DFF_626(CK,g3602,g30428);
  FD1 DFF_627(CK,g5571,g30485);
  FD1 DFF_628(CK,g3578,g30422);
  FD1 DFF_629(CK,g468,g25606);
  FD1 DFF_630(CK,g5448,g25714);
  FD1 DFF_631(CK,g3767,g25680);
  FD1 DFF_632(CK,g5827,g29294);
  FD1 DFF_633(CK,g3582,g30423);
  FD1 DFF_634(CK,g6271,g30529);
  FD1 DFF_635(CK,g4688,g34028);
  FD1 DFF_636(CK,g5774,g25724);
  FD1 DFF_637(CK,g2380,g33587);
  FD1 DFF_638(CK,g5196,g30460);
  FD1 DFF_639(CK,g5396,g31910);
  FD1 DFF_640(CK,g3227,g30401);
  FD1 DFF_641(CK,g2020,g33990);
  FD1 DFF_642(CK,g4000,g3976);
  FD1 DFF_643(CK,g1079,g1075);
  FD1 DFF_644(CK,g6541,g29309);
  FD1 DFF_645(CK,g3203,g30411);
  FD1 DFF_646(CK,g1668,g33546);
  FD1 DFF_647(CK,g4760,g28085);
  FD1 DFF_648(CK,g262,g26904);
  FD1 DFF_649(CK,g1840,g33556);
  FD1 DFF_650(CK,g70,g18093);
  FD1 DFF_651(CK,g5467,g25722);
  FD1 DFF_652(CK,g460,g25605);
  FD1 DFF_653(CK,g6209,g33062);
  FD1 DFF_654(CK,g74,g26893);
  FD1 DFF_655(CK,g5290,g5313);
  FD1 DFF_656(CK,g655,g28050);
  FD1 DFF_657(CK,g3502,g34626);
  FD1 DFF_658(CK,g2204,g33583);
  FD1 DFF_659(CK,g5256,g30472);
  FD1 DFF_660(CK,g4608,g34454);
  FD1 DFF_661(CK,g794,g34850);
  FD1 DFF_662(CK,g4023,g4019);
  FD1 DFF_663(CK,g4423,g4537);
  FD1 DFF_664(CK,g3689,g24272);
  FD1 DFF_665(CK,g5381,g31906);
  FD1 DFF_666(CK,g5685,g5681);
  FD1 DFF_667(CK,g703,g24214);
  FD1 DFF_668(CK,g5421,g25718);
  FD1 DFF_669(CK,g862,g26909);
  FD1 DFF_670(CK,g3247,g30406);
  FD1 DFF_671(CK,g2040,g33569);
  FD1 DFF_672(CK,g4999,g25694);
  FD1 DFF_673(CK,g4146,g34628);
  FD1 DFF_674(CK,g4633,g34458);
  FD1 DFF_675(CK,g1157,g24240);
  FD1 DFF_676(CK,g5723,g31918);
  FD1 DFF_677(CK,g4732,g34634);
  FD1 DFF_678(CK,g5101,g25700);
  FD1 DFF_679(CK,g5817,g29293);
  FD1 DFF_680(CK,g2151,g18421);
  FD1 DFF_681(CK,g2351,g33009);
  FD1 DFF_682(CK,g2648,g33603);
  FD1 DFF_683(CK,g6736,g24355);
  FD1 DFF_684(CK,g4944,g34268);
  FD1 DFF_685(CK,g4072,g25691);
  FD1 DFF_686(CK,g344,g26890);
  FD1 DFF_687(CK,g4443,g4449);
  FD1 DFF_688(CK,g3466,g29264);
  FD1 DFF_689(CK,g4116,g28072);
  FD1 DFF_690(CK,g5041,g31900);
  FD1 DFF_691(CK,g5441,g25712);
  FD1 DFF_692(CK,g4434,g26956);
  FD1 DFF_693(CK,g3827,g29271);
  FD1 DFF_694(CK,g6500,g29304);
  FD1 DFF_695(CK,g5673,g5654);
  FD1 DFF_696(CK,g3133,g29261);
  FD1 DFF_697(CK,g3333,g28063);
  FD1 DFF_698(CK,g979,g1116);
  FD1 DFF_699(CK,g4681,g34027);
  FD1 DFF_700(CK,g298,g33961);
  FD1 DFF_701(CK,g3774,g25672);
  FD1 DFF_702(CK,g2667,g33604);
  FD1 DFF_703(CK,g3396,g33025);
  FD1 DFF_704(CK,g4210,g4207);
  FD1 DFF_705(CK,g1894,g32995);
  FD1 DFF_706(CK,g2988,g34624);
  FD1 DFF_707(CK,g3538,g30415);
  FD1 DFF_708(CK,g301,g33536);
  FD1 DFF_709(CK,g341,g26888);
  FD1 DFF_710(CK,g827,g28055);
  FD1 DFF_711(CK,g1075,g24238);
  FD1 DFF_712(CK,g6077,g31921);
  FD1 DFF_713(CK,g2555,g33600);
  FD1 DFF_714(CK,g5011,g28105);
  FD1 DFF_715(CK,g199,g34721);
  FD1 DFF_716(CK,g6523,g29307);
  FD1 DFF_717(CK,g1526,g30345);
  FD1 DFF_718(CK,g4601,g34453);
  FD1 DFF_719(CK,g854,g32980);
  FD1 DFF_720(CK,g1484,g29238);
  FD1 DFF_721(CK,g4922,g34639);
  FD1 DFF_722(CK,g5080,g25695);
  FD1 DFF_723(CK,g5863,g33057);
  FD1 DFF_724(CK,g4581,g26969);
  FD1 DFF_725(CK,g3021,g31879);
  FD1 DFF_726(CK,g2518,g29253);
  FD1 DFF_727(CK,g2567,g34021);
  FD1 DFF_728(CK,g568,g26895);
  FD1 DFF_729(CK,g3263,g30413);
  FD1 DFF_730(CK,g6613,g30549);
  FD1 DFF_731(CK,g6044,g24347);
  FD1 DFF_732(CK,g6444,g25758);
  FD1 DFF_733(CK,g2965,g34808);
  FD1 DFF_734(CK,g5857,g30501);
  FD1 DFF_735(CK,g1616,g33969);
  FD1 DFF_736(CK,g890,g34440);
  FD1 DFF_737(CK,g5976,g5969);
  FD1 DFF_738(CK,g3562,g30433);
  FD1 DFF_739(CK,g4294,g21900);
  FD1 DFF_740(CK,g1404,g26921);
  FD1 DFF_741(CK,g3723,g31893);
  FD1 DFF_742(CK,g3817,g29270);
  FD1 DFF_743(CK,g93,g34878);
  FD1 DFF_744(CK,g4501,g33038);
  FD1 DFF_745(CK,g287,g31865);
  FD1 DFF_746(CK,g2724,g26926);
  FD1 DFF_747(CK,g4704,g28083);
  FD1 DFF_748(CK,g22,g29209);
  FD1 DFF_749(CK,g2878,g34797);
  FD1 DFF_750(CK,g5220,g30478);
  FD1 DFF_751(CK,g617,g34724);
  FD1 DFF_752(CK,g637,g24212);
  FD1 DFF_753(CK,g316,g26883);
  FD1 DFF_754(CK,g1277,g32985);
  FD1 DFF_755(CK,g6513,g25761);
  FD1 DFF_756(CK,g336,g26886);
  FD1 DFF_757(CK,g2882,g34796);
  FD1 DFF_758(CK,g933,g32982);
  FD1 DFF_759(CK,g1906,g33561);
  FD1 DFF_760(CK,g305,g26880);
  FD1 DFF_761(CK,g8,g34591);
  FD1 DFF_762(CK,g3368,g31884);
  FD1 DFF_763(CK,g2799,g26931);
  FD1 DFF_764(CK,g887,g884);
  FD1 DFF_765(CK,g5327,g5308);
  FD1 DFF_766(CK,g4912,g34641);
  FD1 DFF_767(CK,g4157,g34629);
  FD1 DFF_768(CK,g2541,g33598);
  FD1 DFF_769(CK,g2153,g33576);
  FD1 DFF_770(CK,g550,g34720);
  FD1 DFF_771(CK,g255,g26902);
  FD1 DFF_772(CK,g1945,g29244);
  FD1 DFF_773(CK,g5240,g30468);
  FD1 DFF_774(CK,g1478,g26924);
  FD1 DFF_775(CK,g3080,g25645);
  FD1 DFF_776(CK,g3863,g33031);
  FD1 DFF_777(CK,g1959,g29245);
  FD1 DFF_778(CK,g3480,g29266);
  FD1 DFF_779(CK,g6653,g30559);
  FD1 DFF_780(CK,g6719,g6715);
  FD1 DFF_781(CK,g2864,g34794);
  FD1 DFF_782(CK,g4894,g28087);
  FD1 DFF_783(CK,g5681,g5677);
  FD1 DFF_784(CK,g3857,g30435);
  FD1 DFF_785(CK,g3976,g3969);
  FD1 DFF_786(CK,g499,g25609);
  FD1 DFF_787(CK,g5413,g28095);
  FD1 DFF_788(CK,g1002,g28057);
  FD1 DFF_789(CK,g776,g34439);
  FD1 DFF_790(CK,g28,g34595);
  FD1 DFF_791(CK,g1236,g1233);
  FD1 DFF_792(CK,g4646,g34260);
  FD1 DFF_793(CK,g2476,g33012);
  FD1 DFF_794(CK,g1657,g32989);
  FD1 DFF_795(CK,g2375,g34006);
  FD1 DFF_796(CK,g63,g34847);
  FD1 DFF_797(CK,g6012,g5983);
  FD1 DFF_798(CK,g358,g365);
  FD1 DFF_799(CK,g896,g26910);
  FD1 DFF_800(CK,g967,g21722);
  FD1 DFF_801(CK,g3423,g25658);
  FD1 DFF_802(CK,g283,g28043);
  FD1 DFF_803(CK,g3161,g33021);
  FD1 DFF_804(CK,g2384,g29251);
  FD1 DFF_805(CK,g3361,g25665);
  FD1 DFF_806(CK,g6675,g6697);
  FD1 DFF_807(CK,g4616,g34456);
  FD1 DFF_808(CK,g4561,g26968);
  FD1 DFF_809(CK,g2024,g33991);
  FD1 DFF_810(CK,g3451,g3443);
  FD1 DFF_811(CK,g2795,g26930);
  FD1 DFF_812(CK,g613,g34599);
  FD1 DFF_813(CK,g4527,g28082);
  FD1 DFF_814(CK,g1844,g33557);
  FD1 DFF_815(CK,g5937,g30511);
  FD1 DFF_816(CK,g4546,g33045);
  FD1 DFF_817(CK,g3103,g3096);
  FD1 DFF_818(CK,g2523,g30379);
  FD1 DFF_819(CK,g3303,g24267);
  FD1 DFF_820(CK,g2643,g34020);
  FD1 DFF_821(CK,g6109,g28100);
  FD1 DFF_822(CK,g1489,g24249);
  FD1 DFF_823(CK,g5390,g31908);
  FD1 DFF_824(CK,g194,g25592);
  FD1 DFF_825(CK,g2551,g30382);
  FD1 DFF_826(CK,g5156,g29285);
  FD1 DFF_827(CK,g3072,g25644);
  FD1 DFF_828(CK,g1242,g1227);
  FD1 DFF_829(CK,g47,g34992);
  FD1 DFF_830(CK,g3443,g25662);
  FD1 DFF_831(CK,g4277,g21896);
  FD1 DFF_832(CK,g1955,g33563);
  FD1 DFF_833(CK,g6049,g33622);
  FD1 DFF_834(CK,g3034,g31876);
  FD1 DFF_835(CK,g2273,g33582);
  FD1 DFF_836(CK,g6715,g6711);
  FD1 DFF_837(CK,g4771,g28086);
  FD1 DFF_838(CK,g6098,g25744);
  FD1 DFF_839(CK,g3147,g29262);
  FD1 DFF_840(CK,g3347,g24270);
  FD1 DFF_841(CK,g2269,g33581);
  FD1 DFF_842(CK,g191,g194);
  FD1 DFF_843(CK,g2712,g26937);
  FD1 DFF_844(CK,g626,g34849);
  FD1 DFF_845(CK,g2729,g28060);
  FD1 DFF_846(CK,g5357,g33618);
  FD1 DFF_847(CK,g4991,g34038);
  FD1 DFF_848(CK,g6019,g6000);
  FD1 DFF_849(CK,g4709,g34032);
  FD1 DFF_850(CK,g6419,g31927);
  FD1 DFF_851(CK,g6052,g31919);
  FD1 DFF_852(CK,g2927,g34803);
  FD1 DFF_853(CK,g4340,g34459);
  FD1 DFF_854(CK,g5929,g30509);
  FD1 DFF_855(CK,g4907,g34640);
  FD1 DFF_856(CK,g3317,g3298);
  FD1 DFF_857(CK,g4035,g28069);
  FD1 DFF_858(CK,g2946,g21899);
  FD1 DFF_859(CK,g918,g31868);
  FD1 DFF_860(CK,g4082,g26938);
  FD1 DFF_861(CK,g6486,g25756);
  FD1 DFF_862(CK,g2036,g30363);
  FD1 DFF_863(CK,g577,g30334);
  FD1 DFF_864(CK,g1620,g33970);
  FD1 DFF_865(CK,g2831,g30391);
  FD1 DFF_866(CK,g667,g25615);
  FD1 DFF_867(CK,g930,g33540);
  FD1 DFF_868(CK,g3937,g30445);
  FD1 DFF_869(CK,g5782,g25725);
  FD1 DFF_870(CK,g817,g25617);
  FD1 DFF_871(CK,g1249,g24247);
  FD1 DFF_872(CK,g837,g24215);
  FD1 DFF_873(CK,g3668,g3649);
  FD1 DFF_874(CK,g599,g33964);
  FD1 DFF_875(CK,g5475,g25719);
  FD1 DFF_876(CK,g739,g29228);
  FD1 DFF_877(CK,g5949,g30514);
  FD1 DFF_878(CK,g6682,g33627);
  FD1 DFF_879(CK,g6105,g28101);
  FD1 DFF_880(CK,g904,g24231);
  FD1 DFF_881(CK,g2873,g34615);
  FD1 DFF_882(CK,g1854,g30356);
  FD1 DFF_883(CK,g5084,g25696);
  FD1 DFF_884(CK,g5603,g30493);
  FD1 DFF_885(CK,g4222,g4219);
  FD1 DFF_886(CK,g2495,g33594);
  FD1 DFF_887(CK,g2437,g34009);
  FD1 DFF_888(CK,g2102,g30365);
  FD1 DFF_889(CK,g2208,g33004);
  FD1 DFF_890(CK,g2579,g34018);
  FD1 DFF_891(CK,g4064,g25685);
  FD1 DFF_892(CK,g4899,g34040);
  FD1 DFF_893(CK,g2719,g25639);
  FD1 DFF_894(CK,g4785,g34029);
  FD1 DFF_895(CK,g5583,g30488);
  FD1 DFF_896(CK,g781,g34600);
  FD1 DFF_897(CK,g6173,g29300);
  FD1 DFF_898(CK,g6373,g6369);
  FD1 DFF_899(CK,g2917,g34802);
  FD1 DFF_900(CK,g686,g25614);
  FD1 DFF_901(CK,g1252,g28058);
  FD1 DFF_902(CK,g671,g29225);
  FD1 DFF_903(CK,g2265,g33580);
  FD1 DFF_904(CK,g6283,g30532);
  FD1 DFF_905(CK,g6369,g6365);
  FD1 DFF_906(CK,g5276,g5320);
  FD1 DFF_907(CK,g6459,g25760);
  FD1 DFF_908(CK,g901,g25620);
  FD1 DFF_909(CK,g4194,g4188);
  FD1 DFF_910(CK,g5527,g33054);
  FD1 DFF_911(CK,g4489,g26962);
  FD1 DFF_912(CK,g1974,g33564);
  FD1 DFF_913(CK,g1270,g32984);
  FD1 DFF_914(CK,g4966,g34039);
  FD1 DFF_915(CK,g6415,g31932);
  FD1 DFF_916(CK,g6227,g33065);
  FD1 DFF_917(CK,g3929,g30443);
  FD1 DFF_918(CK,g5503,g29291);
  FD1 DFF_919(CK,g4242,g24279);
  FD1 DFF_920(CK,g5925,g30508);
  FD1 DFF_921(CK,g1124,g29232);
  FD1 DFF_922(CK,g4955,g34269);
  FD1 DFF_923(CK,g5224,g30464);
  FD1 DFF_924(CK,g2012,g33988);
  FD1 DFF_925(CK,g6203,g30522);
  FD1 DFF_926(CK,g5120,g25708);
  FD1 DFF_927(CK,g5320,g5290);
  FD1 DFF_928(CK,g2389,g30374);
  FD1 DFF_929(CK,g4438,g26953);
  FD1 DFF_930(CK,g2429,g34008);
  FD1 DFF_931(CK,g2787,g34444);
  FD1 DFF_932(CK,g1287,g34731);
  FD1 DFF_933(CK,g2675,g33606);
  FD1 DFF_934(CK,g66,g24334);
  FD1 DFF_935(CK,g4836,g34265);
  FD1 DFF_936(CK,g1199,g30340);
  FD1 DFF_937(CK,g1399,g24257);
  FD1 DFF_938(CK,g5547,g30482);
  FD1 DFF_939(CK,g3782,g25673);
  FD1 DFF_940(CK,g6428,g31929);
  FD1 DFF_941(CK,g2138,g34604);
  FD1 DFF_942(CK,g3661,g3632);
  FD1 DFF_943(CK,g2338,g33591);
  FD1 DFF_944(CK,g4229,g4226);
  FD1 DFF_945(CK,g6247,g30525);
  FD1 DFF_946(CK,g2791,g26929);
  FD1 DFF_947(CK,g3949,g30448);
  FD1 DFF_948(CK,g1291,g34602);
  FD1 DFF_949(CK,g5945,g30513);
  FD1 DFF_950(CK,g5244,g30469);
  FD1 DFF_951(CK,g2759,g33608);
  FD1 DFF_952(CK,g6741,g33626);
  FD1 DFF_953(CK,g785,g34725);
  FD1 DFF_954(CK,g1259,g30342);
  FD1 DFF_955(CK,g3484,g29267);
  FD1 DFF_956(CK,g209,g25593);
  FD1 DFF_957(CK,g6609,g30548);
  FD1 DFF_958(CK,g5517,g33052);
  FD1 DFF_959(CK,g2449,g34012);
  FD1 DFF_960(CK,g2575,g34017);
  FD1 DFF_961(CK,g65,g34785);
  FD1 DFF_962(CK,g2715,g24263);
  FD1 DFF_963(CK,g936,g26912);
  FD1 DFF_964(CK,g2098,g30364);
  FD1 DFF_965(CK,g4462,g34254);
  FD1 DFF_966(CK,g604,g34251);
  FD1 DFF_967(CK,g6589,g30560);
  FD1 DFF_968(CK,g1886,g33983);
  FD1 DFF_969(CK,g6466,g25752);
  FD1 DFF_970(CK,g6365,g6346);
  FD1 DFF_971(CK,g6711,g6692);
  FD1 DFF_972(CK,g429,g24204);
  FD1 DFF_973(CK,g1870,g33980);
  FD1 DFF_974(CK,g4249,g34631);
  FD1 DFF_975(CK,g6455,g28103);
  FD1 DFF_976(CK,g3004,g31873);
  FD1 DFF_977(CK,g1825,g29243);
  FD1 DFF_978(CK,g6133,g25740);
  FD1 DFF_979(CK,g1008,g25623);
  FD1 DFF_980(CK,g4392,g26950);
  FD1 DFF_981(CK,g5002,g4999);
  FD1 DFF_982(CK,g3546,g30431);
  FD1 DFF_983(CK,g5236,g30467);
  FD1 DFF_984(CK,g1768,g30353);
  FD1 DFF_985(CK,g4854,g34467);
  FD1 DFF_986(CK,g3925,g30442);
  FD1 DFF_987(CK,g6509,g29305);
  FD1 DFF_988(CK,g732,g25616);
  FD1 DFF_989(CK,g2504,g29252);
  FD1 DFF_990(CK,g1322,g1459);
  FD1 DFF_991(CK,g4520,g6972);
  FD1 DFF_992(CK,g4219,g4216);
  FD1 DFF_993(CK,g2185,g33003);
  FD1 DFF_994(CK,g37,g34613);
  FD1 DFF_995(CK,g4031,g4027);
  FD1 DFF_996(CK,g2070,g33570);
  FD1 DFF_997(CK,g4812,g4809);
  FD1 DFF_998(CK,g6093,g33061);
  FD1 DFF_999(CK,g968,g21723);
  FD1 DFF_1000(CK,g4176,g34734);
  FD1 DFF_1001(CK,g4005,g24275);
  FD1 DFF_1002(CK,g4405,g4408);
  FD1 DFF_1003(CK,g872,g887);
  FD1 DFF_1004(CK,g6181,g29302);
  FD1 DFF_1005(CK,g6381,g24349);
  FD1 DFF_1006(CK,g4765,g34264);
  FD1 DFF_1007(CK,g5563,g30484);
  FD1 DFF_1008(CK,g1395,g25634);
  FD1 DFF_1009(CK,g1913,g33567);
  FD1 DFF_1010(CK,g2331,g33585);
  FD1 DFF_1011(CK,g6263,g30527);
  FD1 DFF_1012(CK,g50,g34995);
  FD1 DFF_1013(CK,g3945,g30447);
  FD1 DFF_1014(CK,g347,g344);
  FD1 DFF_1015(CK,g5731,g31914);
  FD1 DFF_1016(CK,g4473,g34256);
  FD1 DFF_1017(CK,g1266,g25630);
  FD1 DFF_1018(CK,g5489,g29290);
  FD1 DFF_1019(CK,g714,g29227);
  FD1 DFF_1020(CK,g2748,g31872);
  FD1 DFF_1021(CK,g5471,g29287);
  FD1 DFF_1022(CK,g4540,g31897);
  FD1 DFF_1023(CK,g6723,g6719);
  FD1 DFF_1024(CK,g6605,g30562);
  FD1 DFF_1025(CK,g2445,g34011);
  FD1 DFF_1026(CK,g2173,g33996);
  FD1 DFF_1027(CK,g4287,g21898);
  FD1 DFF_1028(CK,g2491,g33014);
  FD1 DFF_1029(CK,g4849,g34465);
  FD1 DFF_1030(CK,g2169,g33995);
  FD1 DFF_1031(CK,g2283,g30372);
  FD1 DFF_1032(CK,g6585,g30545);
  FD1 DFF_1033(CK,g121,g30389);
  FD1 DFF_1034(CK,g2407,g33590);
  FD1 DFF_1035(CK,g2868,g34616);
  FD1 DFF_1036(CK,g2767,g26927);
  FD1 DFF_1037(CK,g1783,g32992);
  FD1 DFF_1038(CK,g3310,g3281);
  FD1 DFF_1039(CK,g1312,g25631);
  FD1 DFF_1040(CK,g5212,g30477);
  FD1 DFF_1041(CK,g4245,g34632);
  FD1 DFF_1042(CK,g645,g28046);
  FD1 DFF_1043(CK,g4291,g4287);
  FD1 DFF_1044(CK,g79,g26896);
  FD1 DFF_1045(CK,g182,g25602);
  FD1 DFF_1046(CK,g1129,g26916);
  FD1 DFF_1047(CK,g2227,g33578);
  FD1 DFF_1048(CK,g6058,g25745);
  FD1 DFF_1049(CK,g4207,g4204);
  FD1 DFF_1050(CK,g2246,g33579);
  FD1 DFF_1051(CK,g1830,g30354);
  FD1 DFF_1052(CK,g3590,g30425);
  FD1 DFF_1053(CK,g392,g24200);
  FD1 DFF_1054(CK,g1592,g33544);
  FD1 DFF_1055(CK,g6505,g25764);
  FD1 DFF_1056(CK,g6411,g31930);
  FD1 DFF_1057(CK,g1221,g24246);
  FD1 DFF_1058(CK,g5921,g30507);
  FD1 DFF_1059(CK,g106,g26889);
  FD1 DFF_1060(CK,g146,g30333);
  FD1 DFF_1061(CK,g218,g215);
  FD1 DFF_1062(CK,g6474,g25753);
  FD1 DFF_1063(CK,g1932,g32998);
  FD1 DFF_1064(CK,g1624,g32987);
  FD1 DFF_1065(CK,g5062,g25702);
  FD1 DFF_1066(CK,g5462,g29286);
  FD1 DFF_1067(CK,g2689,g34606);
  FD1 DFF_1068(CK,g6573,g33070);
  FD1 DFF_1069(CK,g1677,g29240);
  FD1 DFF_1070(CK,g2028,g32999);
  FD1 DFF_1071(CK,g2671,g33605);
  FD1 DFF_1072(CK,g1576,g24255);
  FD1 DFF_1073(CK,g4408,g26945);
  FD1 DFF_1074(CK,g34,g34877);
  FD1 DFF_1075(CK,g1848,g33558);
  FD1 DFF_1076(CK,g3089,g25647);
  FD1 DFF_1077(CK,g3731,g31889);
  FD1 DFF_1078(CK,g86,g25699);
  FD1 DFF_1079(CK,g5485,g29289);
  FD1 DFF_1080(CK,g2741,g30388);
  FD1 DFF_1081(CK,g802,g799);
  FD1 DFF_1082(CK,g2638,g29254);
  FD1 DFF_1083(CK,g4122,g28074);
  FD1 DFF_1084(CK,g4322,g34450);
  FD1 DFF_1085(CK,g5941,g30512);
  FD1 DFF_1086(CK,g2108,g33572);
  FD1 DFF_1087(CK,g6000,g5976);
  FD1 DFF_1088(CK,g25,g15048);
  FD1 DFF_1089(CK,g1644,g33551);
  FD1 DFF_1090(CK,g595,g33538);
  FD1 DFF_1091(CK,g2217,g33005);
  FD1 DFF_1092(CK,g1319,g24248);
  FD1 DFF_1093(CK,g2066,g33002);
  FD1 DFF_1094(CK,g1152,g24234);
  FD1 DFF_1095(CK,g5252,g30471);
  FD1 DFF_1096(CK,g2165,g34000);
  FD1 DFF_1097(CK,g2571,g34016);
  FD1 DFF_1098(CK,g5176,g33048);
  FD1 DFF_1099(CK,g391,g26911);
  FD1 DFF_1100(CK,g5005,g5002);
  FD1 DFF_1101(CK,g2711,g18528);
  FD1 DFF_1102(CK,g6023,g6019);
  FD1 DFF_1103(CK,g1211,g25628);
  FD1 DFF_1104(CK,g2827,g26934);
  FD1 DFF_1105(CK,g6423,g31928);
  FD1 DFF_1106(CK,g875,g869);
  FD1 DFF_1107(CK,g4859,g34468);
  FD1 DFF_1108(CK,g424,g24202);
  FD1 DFF_1109(CK,g1274,g33542);
  FD1 DFF_1110(CK,g1426,g1422);
  FD1 DFF_1111(CK,g85,g34717);
  FD1 DFF_1112(CK,g2803,g34445);
  FD1 DFF_1113(CK,g6451,g28104);
  FD1 DFF_1114(CK,g1821,g33555);
  FD1 DFF_1115(CK,g2509,g34013);
  FD1 DFF_1116(CK,g5073,g28091);
  FD1 DFF_1117(CK,g1280,g26919);
  FD1 DFF_1118(CK,g4815,g4812);
  FD1 DFF_1119(CK,g6346,g6322);
  FD1 DFF_1120(CK,g6633,g30554);
  FD1 DFF_1121(CK,g5124,g29281);
  FD1 DFF_1122(CK,g1083,g1079);
  FD1 DFF_1123(CK,g6303,g30537);
  FD1 DFF_1124(CK,g5069,g28092);
  FD1 DFF_1125(CK,g2994,g34732);
  FD1 DFF_1126(CK,g650,g28049);
  FD1 DFF_1127(CK,g1636,g33545);
  FD1 DFF_1128(CK,g3921,g30441);
  FD1 DFF_1129(CK,g2093,g29247);
  FD1 DFF_1130(CK,g6732,g24354);
  FD1 DFF_1131(CK,g1306,g25636);
  FD1 DFF_1132(CK,g5377,g31911);
  FD1 DFF_1133(CK,g1061,g26914);
  FD1 DFF_1134(CK,g3462,g25670);
  FD1 DFF_1135(CK,g2181,g33998);
  FD1 DFF_1136(CK,g956,g25626);
  FD1 DFF_1137(CK,g1756,g33977);
  FD1 DFF_1138(CK,g5849,g29297);
  FD1 DFF_1139(CK,g4112,g28071);
  FD1 DFF_1140(CK,g2685,g30387);
  FD1 DFF_1141(CK,g2197,g33577);
  FD1 DFF_1142(CK,g6116,g25737);
  FD1 DFF_1143(CK,g2421,g33592);
  FD1 DFF_1144(CK,g1046,g26913);
  FD1 DFF_1145(CK,g482,g28044);
  FD1 DFF_1146(CK,g4401,g26948);
  FD1 DFF_1147(CK,g6434,g31931);
  FD1 DFF_1148(CK,g1514,g30344);
  FD1 DFF_1149(CK,g329,g26885);
  FD1 DFF_1150(CK,g6565,g33069);
  FD1 DFF_1151(CK,g2950,g34621);
  FD1 DFF_1152(CK,g4129,g28075);
  FD1 DFF_1153(CK,g1345,g28059);
  FD1 DFF_1154(CK,g6533,g25762);
  FD1 DFF_1155(CK,g3298,g3274);
  FD1 DFF_1156(CK,g3085,g25646);
  FD1 DFF_1157(CK,g4727,g34633);
  FD1 DFF_1158(CK,g6697,g24352);
  FD1 DFF_1159(CK,g1536,g26925);
  FD1 DFF_1160(CK,g3941,g30446);
  FD1 DFF_1161(CK,g370,g25597);
  FD1 DFF_1162(CK,g5694,g24342);
  FD1 DFF_1163(CK,g1858,g30357);
  FD1 DFF_1164(CK,g446,g26908);
  FD1 DFF_1165(CK,g4932,g21905);
  FD1 DFF_1166(CK,g3219,g30399);
  FD1 DFF_1167(CK,g1811,g29242);
  FD1 DFF_1168(CK,g3431,g25659);
  FD1 DFF_1169(CK,g6601,g30547);
  FD1 DFF_1170(CK,g3376,g31881);
  FD1 DFF_1171(CK,g2441,g34010);
  FD1 DFF_1172(CK,g1874,g33986);
  FD1 DFF_1173(CK,g4349,g34257);
  FD1 DFF_1174(CK,g6581,g30544);
  FD1 DFF_1175(CK,g6597,g30561);
  FD1 DFF_1176(CK,g5008,g5005);
  FD1 DFF_1177(CK,g3610,g30430);
  FD1 DFF_1178(CK,g2890,g34799);
  FD1 DFF_1179(CK,g1978,g33565);
  FD1 DFF_1180(CK,g1612,g33968);
  FD1 DFF_1181(CK,g112,g34879);
  FD1 DFF_1182(CK,g2856,g34793);
  FD1 DFF_1183(CK,g6479,g25754);
  FD1 DFF_1184(CK,g1982,g33566);
  FD1 DFF_1185(CK,g6668,g6661);
  FD1 DFF_1186(CK,g5228,g30465);
  FD1 DFF_1187(CK,g4119,g28073);
  FD1 DFF_1188(CK,g6390,g24351);
  FD1 DFF_1189(CK,g1542,g30346);
  FD1 DFF_1190(CK,g4258,g21893);
  FD1 DFF_1191(CK,g4818,g4815);
  FD1 DFF_1192(CK,g5033,g31904);
  FD1 DFF_1193(CK,g4717,g34635);
  FD1 DFF_1194(CK,g1554,g25637);
  FD1 DFF_1195(CK,g3849,g29274);
  FD1 DFF_1196(CK,g6704,g6675);
  FD1 DFF_1197(CK,g3199,g30396);
  FD1 DFF_1198(CK,g5845,g25735);
  FD1 DFF_1199(CK,g4975,g34037);
  FD1 DFF_1200(CK,g790,g34791);
  FD1 DFF_1201(CK,g5913,g30520);
  FD1 DFF_1202(CK,g1902,g30358);
  FD1 DFF_1203(CK,g6163,g29299);
  FD1 DFF_1204(CK,g4125,g28081);
  FD1 DFF_1205(CK,g4821,g28096);
  FD1 DFF_1206(CK,g4939,g28088);
  FD1 DFF_1207(CK,g1056,g24241);
  FD1 DFF_1208(CK,g3207,g30397);
  FD1 DFF_1209(CK,g4483,g4520);
  FD1 DFF_1210(CK,g3259,g30409);
  FD1 DFF_1211(CK,g5142,g29284);
  FD1 DFF_1212(CK,g5248,g30470);
  FD1 DFF_1213(CK,g2126,g30367);
  FD1 DFF_1214(CK,g3694,g24273);
  FD1 DFF_1215(CK,g5481,g29288);
  FD1 DFF_1216(CK,g1964,g30359);
  FD1 DFF_1217(CK,g5097,g25698);
  FD1 DFF_1218(CK,g3215,g30398);
  FD1 DFF_1219(CK,g4027,g4023);
  FD1 DFF_1220(CK,g111,g34718);
  FD1 DFF_1221(CK,g4427,g26952);
  FD1 DFF_1222(CK,g7,g34590);
  FD1 DFF_1223(CK,g2779,g26928);
  FD1 DFF_1224(CK,g4200,g4197);
  FD1 DFF_1225(CK,g4446,g26954);
  FD1 DFF_1226(CK,g1720,g30351);
  FD1 DFF_1227(CK,g1367,g31871);
  FD1 DFF_1228(CK,g5112,g5105);
  FD1 DFF_1229(CK,g19,g34594);
  FD1 DFF_1230(CK,g4145,g26939);
  FD1 DFF_1231(CK,g2161,g33994);
  FD1 DFF_1232(CK,g376,g25596);
  FD1 DFF_1233(CK,g2361,g33586);
  FD1 DFF_1234(CK,g4191,g21901);
  FD1 DFF_1235(CK,g582,g31866);
  FD1 DFF_1236(CK,g2051,g33000);
  FD1 DFF_1237(CK,g1193,g26918);
  FD1 DFF_1238(CK,g5401,g33051);
  FD1 DFF_1239(CK,g3408,g28065);
  FD1 DFF_1240(CK,g2327,g30373);
  FD1 DFF_1241(CK,g907,g28056);
  FD1 DFF_1242(CK,g947,g34601);
  FD1 DFF_1243(CK,g1834,g30355);
  FD1 DFF_1244(CK,g3594,g30426);
  FD1 DFF_1245(CK,g2999,g34805);
  FD1 DFF_1246(CK,g5727,g31913);
  FD1 DFF_1247(CK,g2303,g34002);
  FD1 DFF_1248(CK,g6661,g6704);
  FD1 DFF_1249(CK,g3065,g25652);
  FD1 DFF_1250(CK,g699,g28053);
  FD1 DFF_1251(CK,g723,g29229);
  FD1 DFF_1252(CK,g5703,g33620);
  FD1 DFF_1253(CK,g546,g34722);
  FD1 DFF_1254(CK,g2472,g33599);
  FD1 DFF_1255(CK,g5953,g30515);
  FD1 DFF_1256(CK,g3096,g25649);
  FD1 DFF_1257(CK,g6439,g33066);
  FD1 DFF_1258(CK,g1740,g33979);
  FD1 DFF_1259(CK,g3550,g30417);
  FD1 DFF_1260(CK,g3845,g25683);
  FD1 DFF_1261(CK,g2116,g33574);
  FD1 DFF_1262(CK,g5677,g5673);
  FD1 DFF_1263(CK,g3195,g30410);
  FD1 DFF_1264(CK,g3913,g30454);
  FD1 DFF_1265(CK,g4537,g34024);
  FD1 DFF_1266(CK,g1687,g33547);
  FD1 DFF_1267(CK,g2681,g30386);
  FD1 DFF_1268(CK,g2533,g33596);
  FD1 DFF_1269(CK,g324,g26887);
  FD1 DFF_1270(CK,g2697,g34607);
  FD1 DFF_1271(CK,g5747,g33056);
  FD1 DFF_1272(CK,g4417,g31895);
  FD1 DFF_1273(CK,g6561,g33068);
  FD1 DFF_1274(CK,g1141,g29233);
  FD1 DFF_1275(CK,g1570,g24258);
  FD1 DFF_1276(CK,g2413,g30376);
  FD1 DFF_1277(CK,g1710,g33549);
  FD1 DFF_1278(CK,g6527,g29308);
  FD1 DFF_1279(CK,g6404,g25759);
  FD1 DFF_1280(CK,g3255,g30408);
  FD1 DFF_1281(CK,g1691,g29241);
  FD1 DFF_1282(CK,g2936,g34620);
  FD1 DFF_1283(CK,g5644,g33621);
  FD1 DFF_1284(CK,g5152,g25707);
  FD1 DFF_1285(CK,g5352,g24339);
  FD1 DFF_1286(CK,g4213,g4185);
  FD1 DFF_1287(CK,g6120,g25738);
  FD1 DFF_1288(CK,g2775,g34443);
  FD1 DFF_1289(CK,g2922,g34619);
  FD1 DFF_1290(CK,g1111,g29234);
  FD1 DFF_1291(CK,g5893,g30503);
  FD1 DFF_1292(CK,g1311,g21724);
  FD1 DFF_1293(CK,g3267,g3310);
  FD1 DFF_1294(CK,g6617,g30550);
  FD1 DFF_1295(CK,g2060,g33001);
  FD1 DFF_1296(CK,g4512,g33040);
  FD1 DFF_1297(CK,g5599,g30492);
  FD1 DFF_1298(CK,g3401,g25664);
  FD1 DFF_1299(CK,g4366,g26944);
  FD1 DFF_1300(CK,g3676,g3672);
  FD1 DFF_1301(CK,g94,g34614);
  FD1 DFF_1302(CK,g3129,g29260);
  FD1 DFF_1303(CK,g3329,g3325);
  FD1 DFF_1304(CK,g5170,g33047);
  FD1 DFF_1305(CK,g4456,g25692);
  FD1 DFF_1306(CK,g5821,g25733);
  FD1 DFF_1307(CK,g6299,g30536);
  FD1 DFF_1308(CK,g1239,g1157);
  FD1 DFF_1309(CK,g3727,g31888);
  FD1 DFF_1310(CK,g2079,g29246);
  FD1 DFF_1311(CK,g4698,g34261);
  FD1 DFF_1312(CK,g3703,g33611);
  FD1 DFF_1313(CK,g1559,g25638);
  FD1 DFF_1314(CK,g943,g34728);
  FD1 DFF_1315(CK,g411,g29222);
  FD1 DFF_1316(CK,g6140,g25742);
  FD1 DFF_1317(CK,g3953,g30449);
  FD1 DFF_1318(CK,g3068,g25643);
  FD1 DFF_1319(CK,g2704,g34608);
  FD1 DFF_1320(CK,g6035,g24345);
  FD1 DFF_1321(CK,g6082,g31922);
  FD1 DFF_1322(CK,g49,g34994);
  FD1 DFF_1323(CK,g1300,g25635);
  FD1 DFF_1324(CK,g4057,g25686);
  FD1 DFF_1325(CK,g5200,g30461);
  FD1 DFF_1326(CK,g4843,g34466);
  FD1 DFF_1327(CK,g5046,g31901);
  FD1 DFF_1328(CK,g2250,g29249);
  FD1 DFF_1329(CK,g319,g26882);
  FD1 DFF_1330(CK,g4549,g33041);
  FD1 DFF_1331(CK,g2453,g33011);
  FD1 DFF_1332(CK,g5841,g25734);
  FD1 DFF_1333(CK,g5763,g28097);
  FD1 DFF_1334(CK,g3747,g33030);
  FD1 DFF_1335(CK,g5637,g5659);
  FD1 DFF_1336(CK,g2912,g34618);
  FD1 DFF_1337(CK,g2357,g33010);
  FD1 DFF_1338(CK,g4232,g4229);
  FD1 DFF_1339(CK,g164,g31864);
  FD1 DFF_1340(CK,g4253,g34630);
  FD1 DFF_1341(CK,g5016,g31898);
  FD1 DFF_1342(CK,g3119,g25653);
  FD1 DFF_1343(CK,g1351,g25632);
  FD1 DFF_1344(CK,g1648,g32988);
  FD1 DFF_1345(CK,g4519,g33616);
  FD1 DFF_1346(CK,g5115,g29280);
  FD1 DFF_1347(CK,g3352,g33609);
  FD1 DFF_1348(CK,g6657,g30563);
  FD1 DFF_1349(CK,g4552,g33044);
  FD1 DFF_1350(CK,g3893,g30437);
  FD1 DFF_1351(CK,g3211,g30412);
  FD1 DFF_1352(CK,g5654,g5630);
  FD1 DFF_1353(CK,g929,g21725);
  FD1 DFF_1354(CK,g3274,g3267);
  FD1 DFF_1355(CK,g5595,g30491);
  FD1 DFF_1356(CK,g3614,g30434);
  FD1 DFF_1357(CK,g2894,g34612);
  FD1 DFF_1358(CK,g3125,g29259);
  FD1 DFF_1359(CK,g3325,g3321);
  FD1 DFF_1360(CK,g3821,g25681);
  FD1 DFF_1361(CK,g4141,g25687);
  FD1 DFF_1362(CK,g4570,g33617);
  FD1 DFF_1363(CK,g5272,g30479);
  FD1 DFF_1364(CK,g2735,g29256);
  FD1 DFF_1365(CK,g728,g28054);
  FD1 DFF_1366(CK,g6295,g30535);
  FD1 DFF_1367(CK,g5417,g28094);
  FD1 DFF_1368(CK,g2661,g30385);
  FD1 DFF_1369(CK,g1988,g30361);
  FD1 DFF_1370(CK,g5128,g25705);
  FD1 DFF_1371(CK,g1548,g24260);
  FD1 DFF_1372(CK,g3106,g29257);
  FD1 DFF_1373(CK,g4659,g34461);
  FD1 DFF_1374(CK,g4358,g34258);
  FD1 DFF_1375(CK,g1792,g32993);
  FD1 DFF_1376(CK,g2084,g33992);
  FD1 DFF_1377(CK,g3061,g28061);
  FD1 DFF_1378(CK,g3187,g30394);
  FD1 DFF_1379(CK,g4311,g34449);
  FD1 DFF_1380(CK,g2583,g34019);
  FD1 DFF_1381(CK,g3003,g21726);
  FD1 DFF_1382(CK,g1094,g29231);
  FD1 DFF_1383(CK,g3841,g25682);
  FD1 DFF_1384(CK,g4284,g21897);
  FD1 DFF_1385(CK,g3763,g28067);
  FD1 DFF_1386(CK,g3191,g30395);
  FD1 DFF_1387(CK,g4239,g21892);
  FD1 DFF_1388(CK,g3391,g31885);
  FD1 DFF_1389(CK,g4180,g4210);
  FD1 DFF_1390(CK,g691,g28048);
  FD1 DFF_1391(CK,g534,g34723);
  FD1 DFF_1392(CK,g5366,g25717);
  FD1 DFF_1393(CK,g385,g25598);
  FD1 DFF_1394(CK,g2004,g33987);
  FD1 DFF_1395(CK,g2527,g30380);
  FD1 DFF_1396(CK,g5456,g5448);
  FD1 DFF_1397(CK,g4420,g26965);
  FD1 DFF_1398(CK,g5148,g25706);
  FD1 DFF_1399(CK,g4507,g30458);
  FD1 DFF_1400(CK,g5348,g24338);
  FD1 DFF_1401(CK,g3223,g30400);
  FD1 DFF_1402(CK,g4931,g21904);
  FD1 DFF_1403(CK,g2970,g34623);
  FD1 DFF_1404(CK,g5698,g24343);
  FD1 DFF_1405(CK,g3416,g25666);
  FD1 DFF_1406(CK,g5260,g30473);
  FD1 DFF_1407(CK,g1521,g24252);
  FD1 DFF_1408(CK,g3522,g33028);
  FD1 DFF_1409(CK,g3115,g29258);
  FD1 DFF_1410(CK,g3251,g30407);
  FD1 DFF_1411(CK,g1,g26958);
  FD1 DFF_1412(CK,g4628,g34457);
  FD1 DFF_1413(CK,g1996,g33568);
  FD1 DFF_1414(CK,g3447,g25663);
  FD1 DFF_1415(CK,g4515,g26964);
  FD1 DFF_1416(CK,g4204,g4200);
  FD1 DFF_1417(CK,g4300,g34735);
  FD1 DFF_1418(CK,g1724,g30352);
  FD1 DFF_1419(CK,g1379,g33543);
  FD1 DFF_1420(CK,g3654,g24271);
  FD1 DFF_1421(CK,g12,g30326);
  FD1 DFF_1422(CK,g1878,g33981);
  FD1 DFF_1423(CK,g5619,g30500);
  FD1 DFF_1424(CK,g71,g34786);
  FD1 DFF_1425(CK,g59,g29277);
  IV  NOT_0(I28349,g28367);
  IV  NOT_1(g19408,g16066);
  IV  NOT_2(I21294,g18274);
  IV  NOT_3(g13297,g10831);
  IV  NOT_4(g19635,g16349);
  IV  NOT_5(g32394,g30601);
  IV  NOT_6(I19778,g17781);
  IV  NOT_7(g9900,g6);
  IV  NOT_8(g11889,g9954);
  IV  NOT_9(g13103,g10905);
  IV  NOT_10(g17470,g14454);
  IV  NOT_11(g23499,g20785);
  IV  NOT_12(g6895,g3288);
  IV  NOT_13(g9797,g5441);
  IV  NOT_14(g31804,g29385);
  IV  NOT_15(g6837,g968);
  IV  NOT_16(I15824,g1116);
  IV  NOT_17(g20066,g17433);
  IV  NOT_18(g33804,g33250);
  IV  NOT_19(g20231,g17821);
  IV  NOT_20(I19786,g17844);
  IV  NOT_21(g24066,g21127);
  IV  NOT_22(g11888,g10160);
  IV  NOT_23(g9510,g5835);
  IV  NOT_24(I22692,g21308);
  IV  NOT_25(g12884,g10392);
  IV  NOT_26(g22494,g19801);
  IV  NOT_27(g9245,I13031);
  IV  NOT_28(g8925,I12910);
  IV  NOT_29(g34248,I32243);
  IV  NOT_30(g10289,g1319);
  IV  NOT_31(g11181,g8134);
  IV  NOT_32(I20116,g15737);
  IV  NOT_33(g7888,g1536);
  IV  NOT_34(g9291,g3021);
  IV  NOT_35(g28559,g27700);
  IV  NOT_36(g21056,g15426);
  IV  NOT_37(I33246,g34970);
  IV  NOT_38(g10288,I13718);
  IV  NOT_39(g8224,g3774);
  IV  NOT_40(g21611,I21210);
  IV  NOT_41(g16718,I17932);
  IV  NOT_42(g21722,I21285);
  IV  NOT_43(I12530,g4815);
  IV  NOT_44(g16521,g13543);
  IV  NOT_45(I22400,g19620);
  IV  NOT_46(g23611,g18833);
  IV  NOT_47(g10571,g10233);
  IV  NOT_48(g17467,g14339);
  IV  NOT_49(g17494,g14339);
  IV  NOT_50(g10308,g4459);
  IV  NOT_51(g27015,g26869);
  IV  NOT_52(g23988,g19277);
  IV  NOT_53(g23924,g18997);
  IV  NOT_54(g12217,I15070);
  IV  NOT_55(g14571,I16688);
  IV  NOT_56(g32318,g31596);
  IV  NOT_57(g32446,g31596);
  IV  NOT_58(g14308,I16471);
  IV  NOT_59(I24041,g22182);
  IV  NOT_60(I14935,g9902);
  IV  NOT_61(g34778,I32976);
  IV  NOT_62(g20511,g17929);
  IV  NOT_63(g26672,g25275);
  IV  NOT_64(g11931,I14749);
  IV  NOT_65(g20763,I20816);
  IV  NOT_66(g23432,g21514);
  IV  NOT_67(I18165,g13177);
  IV  NOT_68(I18523,g14443);
  IV  NOT_69(g21271,I21002);
  IV  NOT_70(I31776,g33204);
  IV  NOT_71(g23271,g20785);
  IV  NOT_72(g22155,g19074);
  IV  NOT_73(I22539,g19606);
  IV  NOT_74(I32231,g34123);
  IV  NOT_75(g34786,I32988);
  IV  NOT_76(g9259,g5176);
  IV  NOT_77(I15190,g6005);
  IV  NOT_78(g17782,I18788);
  IV  NOT_79(g8277,I12483);
  IV  NOT_80(g9819,g92);
  IV  NOT_81(I16969,g13943);
  IV  NOT_82(g32540,g30614);
  IV  NOT_83(g25027,I24191);
  IV  NOT_84(g19711,g17062);
  IV  NOT_85(g22170,g19210);
  IV  NOT_86(g13190,g10939);
  IV  NOT_87(g7297,g6069);
  IV  NOT_88(g17419,g14965);
  IV  NOT_89(g20660,g17873);
  IV  NOT_90(g16861,I18051);
  IV  NOT_91(g21461,g15348);
  IV  NOT_92(g10816,I14054);
  IV  NOT_93(g28713,g27907);
  IV  NOT_94(g15755,g13134);
  IV  NOT_95(g23461,g18833);
  IV  NOT_96(I24237,g23823);
  IV  NOT_97(g34945,g34933);
  IV  NOT_98(g8789,I12779);
  IV  NOT_99(g31833,g29385);
  IV  NOT_100(I18006,g13638);
  IV  NOT_101(I20035,g15706);
  IV  NOT_102(I17207,g13835);
  IV  NOT_103(g30999,g29722);
  IV  NOT_104(g25249,g22228);
  IV  NOT_105(g9488,g1878);
  IV  NOT_106(g19537,g15938);
  IV  NOT_107(g17155,I18205);
  IV  NOT_108(I16855,g10473);
  IV  NOT_109(g15563,I17140);
  IV  NOT_110(g23031,g19801);
  IV  NOT_111(g30090,g29134);
  IV  NOT_112(g30998,g29719);
  IV  NOT_113(g25248,g22228);
  IV  NOT_114(g23650,g20653);
  IV  NOT_115(g7138,g5360);
  IV  NOT_116(g16099,g13437);
  IV  NOT_117(g34998,g34981);
  IV  NOT_118(g23887,g18997);
  IV  NOT_119(g25552,g22594);
  IV  NOT_120(g20916,g18008);
  IV  NOT_121(g27084,g26673);
  IV  NOT_122(g30182,I28419);
  IV  NOT_123(g7963,g4146);
  IV  NOT_124(g10374,g6903);
  IV  NOT_125(I32763,g34511);
  IV  NOT_126(g19606,g17614);
  IV  NOT_127(g19492,g16349);
  IV  NOT_128(g22167,g19074);
  IV  NOT_129(g22194,I21776);
  IV  NOT_130(g7109,g5011);
  IV  NOT_131(g7791,I12199);
  IV  NOT_132(g34672,I32800);
  IV  NOT_133(g16777,I18003);
  IV  NOT_134(g20550,g15864);
  IV  NOT_135(g23529,g20558);
  IV  NOT_136(g6854,g2685);
  IV  NOT_137(g18930,g15789);
  IV  NOT_138(g13024,g11900);
  IV  NOT_139(g32902,g30673);
  IV  NOT_140(g6941,g3990);
  IV  NOT_141(g12110,I14970);
  IV  NOT_142(g32957,g31672);
  IV  NOT_143(g9951,g6133);
  IV  NOT_144(g32377,g30984);
  IV  NOT_145(g12922,g12297);
  IV  NOT_146(g23528,g18833);
  IV  NOT_147(g12321,g9637);
  IV  NOT_148(g28678,g27800);
  IV  NOT_149(g32739,g30735);
  IV  NOT_150(g21393,g17264);
  IV  NOT_151(g23843,g19147);
  IV  NOT_152(g26026,I25105);
  IV  NOT_153(g25081,g22342);
  IV  NOT_154(g20085,g16187);
  IV  NOT_155(g23393,g20739);
  IV  NOT_156(g19750,g16326);
  IV  NOT_157(g30331,I28594);
  IV  NOT_158(g24076,g19984);
  IV  NOT_159(g24085,g20857);
  IV  NOT_160(g17589,g14981);
  IV  NOT_161(g20596,I20690);
  IV  NOT_162(g34932,g34914);
  IV  NOT_163(g23764,g21308);
  IV  NOT_164(g25786,g24518);
  IV  NOT_165(I25869,g25851);
  IV  NOT_166(g32738,g31376);
  IV  NOT_167(g32562,g30673);
  IV  NOT_168(g32645,g30825);
  IV  NOT_169(g14669,g12301);
  IV  NOT_170(g20054,g17328);
  IV  NOT_171(I26337,g26835);
  IV  NOT_172(g24054,g19919);
  IV  NOT_173(I20130,g15748);
  IV  NOT_174(g17588,g14782);
  IV  NOT_175(g17524,g14933);
  IV  NOT_176(I18600,g5335);
  IV  NOT_177(g23869,g19277);
  IV  NOT_178(g32699,g31528);
  IV  NOT_179(g10392,g6989);
  IV  NOT_180(I28576,g28431);
  IV  NOT_181(I28585,g30217);
  IV  NOT_182(I15987,g12381);
  IV  NOT_183(g14668,g12450);
  IV  NOT_184(g25356,g22763);
  IV  NOT_185(g24431,g22722);
  IV  NOT_186(g29725,g28349);
  IV  NOT_187(I15250,g9152);
  IV  NOT_188(g28294,g27295);
  IV  NOT_189(g8945,g608);
  IV  NOT_190(g10489,g9259);
  IV  NOT_191(g11987,I14833);
  IV  NOT_192(g13625,g10971);
  IV  NOT_193(I25161,g24920);
  IV  NOT_194(g17477,g14848);
  IV  NOT_195(g23868,g19277);
  IV  NOT_196(g32698,g30614);
  IV  NOT_197(g31812,g29385);
  IV  NOT_198(g11250,g7502);
  IV  NOT_199(g25380,g23776);
  IV  NOT_200(I32550,g34398);
  IV  NOT_201(g7957,g1252);
  IV  NOT_202(g13250,I15811);
  IV  NOT_203(g20269,g15844);
  IV  NOT_204(g34505,g34409);
  IV  NOT_205(g7049,g5853);
  IV  NOT_206(g20773,I20830);
  IV  NOT_207(g25090,g23630);
  IV  NOT_208(g6958,g4372);
  IV  NOT_209(g20268,g18008);
  IV  NOT_210(g14424,g11136);
  IV  NOT_211(g34717,I32881);
  IV  NOT_212(g12417,g7175);
  IV  NOT_213(g25182,g22763);
  IV  NOT_214(g12936,g12601);
  IV  NOT_215(g20655,I20753);
  IV  NOT_216(g8340,g3050);
  IV  NOT_217(g13943,I16231);
  IV  NOT_218(g21225,g17428);
  IV  NOT_219(g24156,I23312);
  IV  NOT_220(g23259,g21070);
  IV  NOT_221(g24655,g23067);
  IV  NOT_222(I12109,g749);
  IV  NOT_223(I18063,g14357);
  IV  NOT_224(g7715,g1178);
  IV  NOT_225(g29744,g28431);
  IV  NOT_226(g8478,g3103);
  IV  NOT_227(g20180,g17533);
  IV  NOT_228(g17616,g14309);
  IV  NOT_229(g20670,g15426);
  IV  NOT_230(I29447,g30729);
  IV  NOT_231(g10830,g10087);
  IV  NOT_232(I32243,g34134);
  IV  NOT_233(g22305,g19801);
  IV  NOT_234(g24180,I23384);
  IV  NOT_235(g32632,g31070);
  IV  NOT_236(g31795,I29371);
  IV  NOT_237(g9594,g2307);
  IV  NOT_238(g6829,g1319);
  IV  NOT_239(g7498,g6675);
  IV  NOT_240(g23258,g20924);
  IV  NOT_241(g26811,g25206);
  IV  NOT_242(I16590,g11966);
  IV  NOT_243(g10544,I13906);
  IV  NOT_244(g15573,I17154);
  IV  NOT_245(I27492,g27511);
  IV  NOT_246(g9806,g5782);
  IV  NOT_247(g14544,I16663);
  IV  NOT_248(I14653,g9417);
  IV  NOT_249(I33044,g34775);
  IV  NOT_250(I16741,g5677);
  IV  NOT_251(g25513,g23870);
  IV  NOT_252(g32661,g31070);
  IV  NOT_253(g20993,g15615);
  IV  NOT_254(g32547,g30614);
  IV  NOT_255(g32895,g30673);
  IV  NOT_256(g8876,I12855);
  IV  NOT_257(g24839,g23436);
  IV  NOT_258(g23244,I22343);
  IV  NOT_259(g24993,g22384);
  IV  NOT_260(g22177,g19074);
  IV  NOT_261(g16162,g13437);
  IV  NOT_262(g11855,I14671);
  IV  NOT_263(g20667,g15224);
  IV  NOT_264(g17466,g12983);
  IV  NOT_265(g9887,g5802);
  IV  NOT_266(g6974,I11746);
  IV  NOT_267(g24667,g23112);
  IV  NOT_268(g9934,g5849);
  IV  NOT_269(g21069,g15277);
  IV  NOT_270(g25505,g22228);
  IV  NOT_271(g34433,I32470);
  IV  NOT_272(g34387,g34188);
  IV  NOT_273(g10042,g2671);
  IV  NOT_274(g24131,g21209);
  IV  NOT_275(g32481,g31194);
  IV  NOT_276(g14705,I16803);
  IV  NOT_277(I13321,g6486);
  IV  NOT_278(g18975,g15938);
  IV  NOT_279(g19553,g16782);
  IV  NOT_280(g19862,I20233);
  IV  NOT_281(g30097,g29118);
  IV  NOT_282(g8915,I12884);
  IV  NOT_283(g16629,g13990);
  IV  NOT_284(I16150,g10430);
  IV  NOT_285(g21657,g17657);
  IV  NOT_286(g16472,g14098);
  IV  NOT_287(I20781,g17155);
  IV  NOT_288(g21068,g15277);
  IV  NOT_289(g14255,g12381);
  IV  NOT_290(I21477,g18695);
  IV  NOT_291(g14189,I16391);
  IV  NOT_292(g32551,g30735);
  IV  NOT_293(g32572,g30735);
  IV  NOT_294(g23375,g20924);
  IV  NOT_295(I24781,g24264);
  IV  NOT_296(I33146,g34903);
  IV  NOT_297(g7162,g4521);
  IV  NOT_298(g25212,g22763);
  IV  NOT_299(g7268,g1636);
  IV  NOT_300(I11740,g4519);
  IV  NOT_301(g7362,g1906);
  IV  NOT_302(g12909,g10412);
  IV  NOT_303(g9433,g5148);
  IV  NOT_304(g26850,I25576);
  IV  NOT_305(g12543,g9417);
  IV  NOT_306(g17642,g14691);
  IV  NOT_307(g20502,g15373);
  IV  NOT_308(g10678,I13990);
  IV  NOT_309(I22725,g21250);
  IV  NOT_310(I13740,g85);
  IV  NOT_311(g23879,g19210);
  IV  NOT_312(g20557,I20647);
  IV  NOT_313(g23970,g19277);
  IV  NOT_314(g34343,g34089);
  IV  NOT_315(g20210,g16897);
  IV  NOT_316(I22114,g19935);
  IV  NOT_317(g12908,g10414);
  IV  NOT_318(g20618,g15277);
  IV  NOT_319(g11867,I14679);
  IV  NOT_320(g11894,I14702);
  IV  NOT_321(I11685,g117);
  IV  NOT_322(g8310,g2051);
  IV  NOT_323(g23878,g19147);
  IV  NOT_324(g21337,g15758);
  IV  NOT_325(g20443,g15171);
  IV  NOT_326(g10383,g6978);
  IV  NOT_327(g23337,g20924);
  IV  NOT_328(g19757,g17224);
  IV  NOT_329(g9496,g3303);
  IV  NOT_330(g14383,I16535);
  IV  NOT_331(g17733,g14238);
  IV  NOT_332(I16526,g10430);
  IV  NOT_333(g8663,g3343);
  IV  NOT_334(g10030,g116);
  IV  NOT_335(g23886,g21468);
  IV  NOT_336(I18614,g6315);
  IV  NOT_337(g32490,g30673);
  IV  NOT_338(g10093,g5703);
  IV  NOT_339(g18884,g15938);
  IV  NOT_340(g27242,g26183);
  IV  NOT_341(I14576,g8791);
  IV  NOT_342(g11714,g8107);
  IV  NOT_343(g22166,g18997);
  IV  NOT_344(g11450,I14455);
  IV  NOT_345(I17114,g14358);
  IV  NOT_346(I27192,g27662);
  IV  NOT_347(g23792,g19074);
  IV  NOT_348(g23967,g19210);
  IV  NOT_349(g23994,g19277);
  IV  NOT_350(g32784,g31672);
  IV  NOT_351(g9891,g6173);
  IV  NOT_352(I18320,g13605);
  IV  NOT_353(g28037,g26365);
  IV  NOT_354(g8002,g1389);
  IV  NOT_355(g9337,g1608);
  IV  NOT_356(g9913,g2403);
  IV  NOT_357(g32956,g30825);
  IV  NOT_358(I21285,g18215);
  IV  NOT_359(g11819,g7717);
  IV  NOT_360(g11910,g10185);
  IV  NOT_361(g14065,g11048);
  IV  NOT_362(g7086,g4826);
  IV  NOT_363(g13707,g11360);
  IV  NOT_364(g31829,g29385);
  IV  NOT_365(g32889,g31376);
  IV  NOT_366(g11202,I14267);
  IV  NOT_367(g8236,g4812);
  IV  NOT_368(g33920,I31786);
  IV  NOT_369(I21254,g16540);
  IV  NOT_370(g24039,g21256);
  IV  NOT_371(g25620,I24759);
  IV  NOT_372(g21425,g15509);
  IV  NOT_373(g29221,I27579);
  IV  NOT_374(I17744,g14912);
  IV  NOT_375(g23459,g21611);
  IV  NOT_376(I16917,g10582);
  IV  NOT_377(g20038,g17328);
  IV  NOT_378(g23425,g20751);
  IV  NOT_379(g31828,g29385);
  IV  NOT_380(g32888,g30673);
  IV  NOT_381(I15070,g10108);
  IV  NOT_382(g25097,g22342);
  IV  NOT_383(g32824,g31376);
  IV  NOT_384(g10219,g2697);
  IV  NOT_385(g13055,I15682);
  IV  NOT_386(g9807,g5712);
  IV  NOT_387(I30901,g32407);
  IV  NOT_388(g19673,g16931);
  IV  NOT_389(g24038,g21193);
  IV  NOT_390(g14219,g12381);
  IV  NOT_391(g19397,g16449);
  IV  NOT_392(g21458,g15758);
  IV  NOT_393(g6849,g2551);
  IV  NOT_394(I15590,g11988);
  IV  NOT_395(g28155,I26664);
  IV  NOT_396(I13762,g6755);
  IV  NOT_397(g13070,g11984);
  IV  NOT_398(g23458,I22583);
  IV  NOT_399(g32671,g31528);
  IV  NOT_400(I21036,g17221);
  IV  NOT_401(g34229,g33936);
  IV  NOT_402(g10218,g2527);
  IV  NOT_403(I18034,g13680);
  IV  NOT_404(g16172,g13584);
  IV  NOT_405(g20601,g17433);
  IV  NOT_406(g21010,g15634);
  IV  NOT_407(g11986,I14830);
  IV  NOT_408(g7470,g5623);
  IV  NOT_409(I12483,g3096);
  IV  NOT_410(g17476,g14665);
  IV  NOT_411(g17485,I18408);
  IV  NOT_412(I16077,g10430);
  IV  NOT_413(I14745,g10029);
  IV  NOT_414(g11741,g10033);
  IV  NOT_415(g22907,g20453);
  IV  NOT_416(g23545,g21562);
  IV  NOT_417(g23444,I22561);
  IV  NOT_418(g25369,g22228);
  IV  NOT_419(g32931,g30937);
  IV  NOT_420(g33682,I31515);
  IV  NOT_421(g6900,g3440);
  IV  NOT_422(g19634,g16349);
  IV  NOT_423(g19872,g17015);
  IV  NOT_424(g34716,I32878);
  IV  NOT_425(I20542,g16508);
  IV  NOT_426(I25598,g25424);
  IV  NOT_427(g8928,g4340);
  IV  NOT_428(g29812,g28381);
  IV  NOT_429(I28241,g28709);
  IV  NOT_430(g12841,g10357);
  IV  NOT_431(g22594,I21934);
  IV  NOT_432(I16688,g10981);
  IV  NOT_433(g9815,g6098);
  IV  NOT_434(g8064,g3376);
  IV  NOT_435(I18408,g13017);
  IV  NOT_436(I20913,g16964);
  IV  NOT_437(g23086,g20283);
  IV  NOT_438(I32815,g34470);
  IV  NOT_439(g30310,g28830);
  IV  NOT_440(g8899,g807);
  IV  NOT_441(g11735,g8534);
  IV  NOT_442(g29371,I27735);
  IV  NOT_443(I11908,g4449);
  IV  NOT_444(g9692,g1756);
  IV  NOT_445(g13877,g11350);
  IV  NOT_446(I32601,g34319);
  IV  NOT_447(g8785,I12767);
  IV  NOT_448(g24169,I23351);
  IV  NOT_449(g24791,g23850);
  IV  NOT_450(g9497,I13166);
  IV  NOT_451(I16102,g10430);
  IV  NOT_452(g26681,g25396);
  IV  NOT_453(g20168,g17533);
  IV  NOT_454(g9154,I12994);
  IV  NOT_455(g25133,g23733);
  IV  NOT_456(g34925,I33167);
  IV  NOT_457(I26309,g26825);
  IV  NOT_458(g9354,g2719);
  IV  NOT_459(g27014,g25888);
  IV  NOT_460(I27564,g28166);
  IV  NOT_461(g24168,I23348);
  IV  NOT_462(g23322,I22425);
  IV  NOT_463(g32546,g31170);
  IV  NOT_464(g9960,g6474);
  IV  NOT_465(g22519,g19801);
  IV  NOT_466(g22176,g18997);
  IV  NOT_467(g14201,I16401);
  IV  NOT_468(g26802,I25514);
  IV  NOT_469(g28119,g27008);
  IV  NOT_470(g12835,g10352);
  IV  NOT_471(g7635,g1002);
  IV  NOT_472(g14277,I16455);
  IV  NOT_473(g20666,g15224);
  IV  NOT_474(g13018,I15636);
  IV  NOT_475(I16231,g10520);
  IV  NOT_476(g32024,I29582);
  IV  NOT_477(g25228,g23828);
  IV  NOT_478(I19802,g15727);
  IV  NOT_479(g19574,g16826);
  IV  NOT_480(g7766,I12189);
  IV  NOT_481(g19452,g16326);
  IV  NOT_482(g6819,g1046);
  IV  NOT_483(g16540,I17744);
  IV  NOT_484(I19857,g16640);
  IV  NOT_485(g22154,g19074);
  IV  NOT_486(g7087,g6336);
  IV  NOT_487(I33297,g35000);
  IV  NOT_488(g25011,g22763);
  IV  NOT_489(g32860,g30673);
  IV  NOT_490(I18891,g16676);
  IV  NOT_491(g7487,g1259);
  IV  NOT_492(I33103,g34846);
  IV  NOT_493(g8237,g255);
  IV  NOT_494(g18953,g16077);
  IV  NOT_495(I14761,g7753);
  IV  NOT_496(g19912,g17328);
  IV  NOT_497(g17519,I18460);
  IV  NOT_498(g21561,g15595);
  IV  NOT_499(I12183,g2719);
  IV  NOT_500(g21656,g17700);
  IV  NOT_501(g6923,g3791);
  IV  NOT_502(g26765,g25309);
  IV  NOT_503(I25680,g25641);
  IV  NOT_504(g22935,g20283);
  IV  NOT_505(g17092,g14011);
  IV  NOT_506(g34944,g34932);
  IV  NOT_507(g10037,g1848);
  IV  NOT_508(I32791,g34578);
  IV  NOT_509(g32497,g30673);
  IV  NOT_510(g21295,g17533);
  IV  NOT_511(g23353,g20924);
  IV  NOT_512(g29507,g28353);
  IV  NOT_513(I32884,g34690);
  IV  NOT_514(g8844,I12826);
  IV  NOT_515(g11402,g7594);
  IV  NOT_516(g17518,g14918);
  IV  NOT_517(g26549,I25391);
  IV  NOT_518(g17154,g14348);
  IV  NOT_519(g22883,g20391);
  IV  NOT_520(g20556,g15483);
  IV  NOT_521(g23823,I22989);
  IV  NOT_522(g17637,g12933);
  IV  NOT_523(g20580,g17328);
  IV  NOT_524(g26548,g25255);
  IV  NOT_525(g10419,g8821);
  IV  NOT_526(g11866,g9883);
  IV  NOT_527(g11917,I14727);
  IV  NOT_528(g32700,g31579);
  IV  NOT_529(I26687,g27880);
  IV  NOT_530(g32659,g30735);
  IV  NOT_531(g21336,g17367);
  IV  NOT_532(g32625,g31070);
  IV  NOT_533(g10352,g6804);
  IV  NOT_534(g23336,g20924);
  IV  NOT_535(I32479,g34302);
  IV  NOT_536(g19592,I20035);
  IV  NOT_537(g34429,I32458);
  IV  NOT_538(g10155,g2643);
  IV  NOT_539(g10418,g8818);
  IV  NOT_540(g12041,I14905);
  IV  NOT_541(g32658,g31579);
  IV  NOT_542(g19780,g16449);
  IV  NOT_543(g16739,g13223);
  IV  NOT_544(g12430,I15250);
  IV  NOT_545(I16660,g10981);
  IV  NOT_546(g34428,I32455);
  IV  NOT_547(I21074,g17766);
  IV  NOT_548(g23966,g19210);
  IV  NOT_549(g22215,g19277);
  IV  NOT_550(g28036,g26365);
  IV  NOT_551(g27237,g26162);
  IV  NOT_552(g32943,g31710);
  IV  NOT_553(g20110,g16897);
  IV  NOT_554(g11706,I14579);
  IV  NOT_555(g24084,g20720);
  IV  NOT_556(g16738,I17956);
  IV  NOT_557(g9761,g2445);
  IV  NOT_558(g13706,g11280);
  IV  NOT_559(g16645,g13756);
  IV  NOT_560(g12465,g7192);
  IV  NOT_561(I11992,g763);
  IV  NOT_562(g24110,g21209);
  IV  NOT_563(g20922,I20891);
  IV  NOT_564(g27983,g26725);
  IV  NOT_565(g20321,g17821);
  IV  NOT_566(g23017,g20453);
  IV  NOT_567(g32644,g30735);
  IV  NOT_568(g33648,I31482);
  IV  NOT_569(I21238,g16540);
  IV  NOT_570(g34690,I32840);
  IV  NOT_571(g6870,g3089);
  IV  NOT_572(g9828,g2024);
  IV  NOT_573(g20179,g17249);
  IV  NOT_574(g34549,I32617);
  IV  NOT_575(g8948,g785);
  IV  NOT_576(g20531,g15907);
  IV  NOT_577(g12983,I15600);
  IV  NOT_578(g24179,I23381);
  IV  NOT_579(g16290,g13260);
  IV  NOT_580(g32969,g30735);
  IV  NOT_581(g13280,I15846);
  IV  NOT_582(g6825,g979);
  IV  NOT_583(g33755,I31610);
  IV  NOT_584(g17501,I18434);
  IV  NOT_585(g7369,g1996);
  IV  NOT_586(g27142,g26105);
  IV  NOT_587(g8955,g1418);
  IV  NOT_588(g20178,g16971);
  IV  NOT_589(g10194,g6741);
  IV  NOT_590(g19396,g16431);
  IV  NOT_591(g17577,I18504);
  IV  NOT_592(g13624,g10951);
  IV  NOT_593(I14241,g8356);
  IV  NOT_594(I21941,g18918);
  IV  NOT_595(g24178,I23378);
  IV  NOT_596(g14167,I16371);
  IV  NOT_597(g32968,g31376);
  IV  NOT_598(g19731,g17093);
  IV  NOT_599(g29920,g28824);
  IV  NOT_600(g34504,g34408);
  IV  NOT_601(g29358,I27718);
  IV  NOT_602(g7868,g1099);
  IV  NOT_603(I15102,g5313);
  IV  NOT_604(I26195,g26260);
  IV  NOT_605(I11835,g101);
  IV  NOT_606(I20891,g17700);
  IV  NOT_607(g9746,I13326);
  IV  NOT_608(g20373,g17929);
  IV  NOT_609(g32855,g30825);
  IV  NOT_610(g23289,g20924);
  IV  NOT_611(g24685,g23139);
  IV  NOT_612(g24373,g22908);
  IV  NOT_613(I33024,g34783);
  IV  NOT_614(g8150,g2185);
  IV  NOT_615(g10401,g7041);
  IV  NOT_616(g22906,g20453);
  IV  NOT_617(g20654,I20750);
  IV  NOT_618(I16596,g12640);
  IV  NOT_619(g34317,g34115);
  IV  NOT_620(g8350,g4646);
  IV  NOT_621(g18908,g16100);
  IV  NOT_622(g32870,g31021);
  IV  NOT_623(g7535,g1500);
  IV  NOT_624(g32527,g30673);
  IV  NOT_625(I13007,g65);
  IV  NOT_626(g8038,I12360);
  IV  NOT_627(g10119,g2841);
  IV  NOT_628(I24474,g22546);
  IV  NOT_629(g16632,g14454);
  IV  NOT_630(g21308,g17485);
  IV  NOT_631(g8438,g3100);
  IV  NOT_632(g23571,g18833);
  IV  NOT_633(g28693,g27837);
  IV  NOT_634(g23308,g21024);
  IV  NOT_635(g31794,I29368);
  IV  NOT_636(g6972,I11740);
  IV  NOT_637(g31845,g29385);
  IV  NOT_638(g8009,g3106);
  IV  NOT_639(I31497,g33187);
  IV  NOT_640(g7261,g4449);
  IV  NOT_641(g24417,g22171);
  IV  NOT_642(g33845,I31694);
  IV  NOT_643(g10118,g2541);
  IV  NOT_644(I19775,g17780);
  IV  NOT_645(g9932,g5805);
  IV  NOT_646(g28166,I26687);
  IV  NOT_647(g28009,I26516);
  IV  NOT_648(g16661,g14454);
  IV  NOT_649(I17507,g13416);
  IV  NOT_650(g25549,g22763);
  IV  NOT_651(g13876,g11432);
  IV  NOT_652(g13885,g10862);
  IV  NOT_653(g32503,g31194);
  IV  NOT_654(g23495,I22622);
  IV  NOT_655(I31659,g33219);
  IV  NOT_656(g14749,I16829);
  IV  NOT_657(g32867,g30673);
  IV  NOT_658(g32894,g30614);
  IV  NOT_659(I31625,g33197);
  IV  NOT_660(g14616,I16733);
  IV  NOT_661(g34245,I32234);
  IV  NOT_662(I32953,g34656);
  IV  NOT_663(g8836,g736);
  IV  NOT_664(g30299,g28765);
  IV  NOT_665(g6887,g3333);
  IV  NOT_666(g23816,g21308);
  IV  NOT_667(g25548,g22550);
  IV  NOT_668(g34323,g34105);
  IV  NOT_669(g34299,g34080);
  IV  NOT_670(I32654,g34378);
  IV  NOT_671(g22139,I21722);
  IV  NOT_672(g8918,I12893);
  IV  NOT_673(g24964,I24128);
  IV  NOT_674(g7246,g4446);
  IV  NOT_675(I11746,g4570);
  IV  NOT_676(g26856,I25586);
  IV  NOT_677(g13763,g10971);
  IV  NOT_678(g14276,I16452);
  IV  NOT_679(g31521,I29182);
  IV  NOT_680(I32800,g34582);
  IV  NOT_681(g32581,g31070);
  IV  NOT_682(g32714,g31528);
  IV  NOT_683(g32450,g31591);
  IV  NOT_684(g10053,g6381);
  IV  NOT_685(g23985,g19210);
  IV  NOT_686(g22138,g21370);
  IV  NOT_687(g15739,g13284);
  IV  NOT_688(I26705,g27967);
  IV  NOT_689(g34775,I32967);
  IV  NOT_690(I20750,g16677);
  IV  NOT_691(g20587,g15373);
  IV  NOT_692(g32707,g31579);
  IV  NOT_693(g32819,g30825);
  IV  NOT_694(g9576,g6565);
  IV  NOT_695(g31832,g29385);
  IV  NOT_696(I20982,g16300);
  IV  NOT_697(g23954,I23099);
  IV  NOT_698(g24587,g23112);
  IV  NOT_699(g8229,g3881);
  IV  NOT_700(g9716,g5057);
  IV  NOT_701(I22788,g18940);
  IV  NOT_702(I26679,g27773);
  IV  NOT_703(g12863,g10371);
  IV  NOT_704(g8993,g385);
  IV  NOT_705(g15562,g14943);
  IV  NOT_706(g32818,g30735);
  IV  NOT_707(g10036,g1816);
  IV  NOT_708(g32496,g30614);
  IV  NOT_709(g19787,g17096);
  IV  NOT_710(g16127,g13437);
  IV  NOT_711(g8822,g4975);
  IV  NOT_712(g10177,g1834);
  IV  NOT_713(g20909,g17955);
  IV  NOT_714(g20543,g17955);
  IV  NOT_715(I13684,g128);
  IV  NOT_716(g31861,I29441);
  IV  NOT_717(g9848,g4462);
  IV  NOT_718(g21669,I21230);
  IV  NOT_719(g19357,I19837);
  IV  NOT_720(g17415,g14797);
  IV  NOT_721(g6845,g2126);
  IV  NOT_722(g7502,I11992);
  IV  NOT_723(I15550,g10430);
  IV  NOT_724(g32590,g31154);
  IV  NOT_725(g9699,g2311);
  IV  NOT_726(g9747,I13329);
  IV  NOT_727(g24117,g21209);
  IV  NOT_728(g24000,g19277);
  IV  NOT_729(I33197,g34930);
  IV  NOT_730(g23260,g21070);
  IV  NOT_731(g19743,g17125);
  IV  NOT_732(I14584,g9766);
  IV  NOT_733(g33926,I31796);
  IV  NOT_734(g25245,g22763);
  IV  NOT_735(g34697,g34545);
  IV  NOT_736(g26831,g24836);
  IV  NOT_737(g20569,g15277);
  IV  NOT_738(I20840,g17727);
  IV  NOT_739(g34995,I33285);
  IV  NOT_740(g23842,g19147);
  IV  NOT_741(g32741,g31710);
  IV  NOT_742(g13314,g10893);
  IV  NOT_743(I23348,g23384);
  IV  NOT_744(g25299,g22763);
  IV  NOT_745(g32384,g31666);
  IV  NOT_746(I19831,g16533);
  IV  NOT_747(g33388,g32382);
  IV  NOT_748(I18252,g13177);
  IV  NOT_749(I16502,g10430);
  IV  NOT_750(g20568,g15509);
  IV  NOT_751(g23489,g21468);
  IV  NOT_752(g25533,g22550);
  IV  NOT_753(g13085,I15717);
  IV  NOT_754(g19769,g16987);
  IV  NOT_755(g24568,g22942);
  IV  NOT_756(g20242,g16308);
  IV  NOT_757(g25298,g23760);
  IV  NOT_758(g11721,g10074);
  IV  NOT_759(g7689,I12159);
  IV  NOT_760(g29927,g28861);
  IV  NOT_761(I17121,g14366);
  IV  NOT_762(g34512,g34420);
  IV  NOT_763(g21424,g15426);
  IV  NOT_764(g23559,g21070);
  IV  NOT_765(g13596,g10971);
  IV  NOT_766(g23525,g21562);
  IV  NOT_767(g23488,g21468);
  IV  NOT_768(g28675,g27779);
  IV  NOT_769(g23016,g20453);
  IV  NOT_770(I32909,g34712);
  IV  NOT_771(g7216,g822);
  IV  NOT_772(g11431,g7618);
  IV  NOT_773(g12952,I15572);
  IV  NOT_774(g23558,g20924);
  IV  NOT_775(g13431,I15932);
  IV  NOT_776(g32801,g30937);
  IV  NOT_777(g14630,g12402);
  IV  NOT_778(g32735,g31021);
  IV  NOT_779(g24123,g21143);
  IV  NOT_780(g32877,g30825);
  IV  NOT_781(g7028,I11785);
  IV  NOT_782(I30686,g32381);
  IV  NOT_783(g8895,g599);
  IV  NOT_784(g10166,g6040);
  IV  NOT_785(g17576,g14953);
  IV  NOT_786(g17585,g14974);
  IV  NOT_787(g20772,g15171);
  IV  NOT_788(g9644,g2016);
  IV  NOT_789(g22200,g19277);
  IV  NOT_790(g23893,g19074);
  IV  NOT_791(I15773,g10430);
  IV  NOT_792(g11269,g7516);
  IV  NOT_793(I15942,g12381);
  IV  NOT_794(g14166,g11048);
  IV  NOT_795(g8620,g3065);
  IV  NOT_796(g19881,g15915);
  IV  NOT_797(g8462,g1183);
  IV  NOT_798(g25232,g22228);
  IV  NOT_799(g29491,I27777);
  IV  NOT_800(g7247,g5377);
  IV  NOT_801(g20639,g15224);
  IV  NOT_802(I17173,g13716);
  IV  NOT_803(g16931,I18101);
  IV  NOT_804(I16468,g12760);
  IV  NOT_805(g23544,g21562);
  IV  NOT_806(g23865,g21308);
  IV  NOT_807(I12046,g613);
  IV  NOT_808(g32695,g30735);
  IV  NOT_809(I31581,g33164);
  IV  NOT_810(g11268,g7515);
  IV  NOT_811(g20230,I20499);
  IV  NOT_812(g12790,g7097);
  IV  NOT_813(g17609,g14817);
  IV  NOT_814(g29755,I28002);
  IV  NOT_815(g7564,g336);
  IV  NOT_816(g9152,g2834);
  IV  NOT_817(g20638,g15224);
  IV  NOT_818(I18509,g5623);
  IV  NOT_819(g9818,g6490);
  IV  NOT_820(g13655,g10573);
  IV  NOT_821(g34316,g34093);
  IV  NOT_822(g17200,I18238);
  IV  NOT_823(g32526,g30614);
  IV  NOT_824(g20265,g17821);
  IV  NOT_825(g29981,g28942);
  IV  NOT_826(g6815,g929);
  IV  NOT_827(I12787,g4311);
  IV  NOT_828(g12873,g10380);
  IV  NOT_829(I22028,g20204);
  IV  NOT_830(I29211,g30298);
  IV  NOT_831(g8788,I12776);
  IV  NOT_832(I18872,g13745);
  IV  NOT_833(I23333,g22683);
  IV  NOT_834(g30989,g29672);
  IV  NOT_835(g33766,I31619);
  IV  NOT_836(g19662,g17432);
  IV  NOT_837(g21610,g15615);
  IV  NOT_838(g14454,I16613);
  IV  NOT_839(g23610,g18833);
  IV  NOT_840(g10570,g9021);
  IV  NOT_841(g34989,I33267);
  IV  NOT_842(g8249,g1917);
  IV  NOT_843(g20391,I20562);
  IV  NOT_844(g32457,g30735);
  IV  NOT_845(g21189,g15634);
  IV  NOT_846(g24992,g22417);
  IV  NOT_847(I33070,g34810);
  IV  NOT_848(g20510,g17226);
  IV  NOT_849(g23189,g20060);
  IV  NOT_850(g11930,g9281);
  IV  NOT_851(g12422,I15238);
  IV  NOT_852(g26736,g25349);
  IV  NOT_853(g9186,I13010);
  IV  NOT_854(g17745,g14978);
  IV  NOT_855(g34988,I33264);
  IV  NOT_856(g22973,g20330);
  IV  NOT_857(g34924,I33164);
  IV  NOT_858(g6960,g1);
  IV  NOT_859(g9386,g5727);
  IV  NOT_860(I15667,g12143);
  IV  NOT_861(I32639,g34345);
  IV  NOT_862(g21270,I20999);
  IV  NOT_863(g32866,g30614);
  IV  NOT_864(g32917,g30937);
  IV  NOT_865(g23270,g20785);
  IV  NOT_866(g19482,g16349);
  IV  NOT_867(g21678,g16540);
  IV  NOT_868(g17813,I18813);
  IV  NOT_869(g12834,g10349);
  IV  NOT_870(g20579,g17249);
  IV  NOT_871(g34432,I32467);
  IV  NOT_872(g7308,g1668);
  IV  NOT_873(g11965,I14797);
  IV  NOT_874(g8085,I12382);
  IV  NOT_875(g9599,g3310);
  IV  NOT_876(g10074,g718);
  IV  NOT_877(g19710,g17059);
  IV  NOT_878(g18983,g16077);
  IV  NOT_879(g24579,g23067);
  IV  NOT_880(g34271,g34160);
  IV  NOT_881(g19552,g16856);
  IV  NOT_882(g21460,g15628);
  IV  NOT_883(g21686,g16540);
  IV  NOT_884(g9274,g5857);
  IV  NOT_885(g20578,g15563);
  IV  NOT_886(g26843,I25567);
  IV  NOT_887(g23460,g21611);
  IV  NOT_888(g23939,g19074);
  IV  NOT_889(g21383,g17367);
  IV  NOT_890(g19779,g16431);
  IV  NOT_891(I19843,g16594);
  IV  NOT_892(g9614,g5128);
  IV  NOT_893(I33067,g34812);
  IV  NOT_894(g17674,I18647);
  IV  NOT_895(g12021,g9543);
  IV  NOT_896(g14238,g10823);
  IV  NOT_897(g20586,g15171);
  IV  NOT_898(g23030,g20453);
  IV  NOT_899(g32706,g30673);
  IV  NOT_900(g23938,g18997);
  IV  NOT_901(g32597,g31154);
  IV  NOT_902(I18574,g13075);
  IV  NOT_903(g25316,g22763);
  IV  NOT_904(g8854,g613);
  IV  NOT_905(g21267,g15680);
  IV  NOT_906(g24586,g23067);
  IV  NOT_907(I32391,g34153);
  IV  NOT_908(g23267,g20097);
  IV  NOT_909(g9821,g115);
  IV  NOT_910(I13236,g5452);
  IV  NOT_911(I18205,g14563);
  IV  NOT_912(g34145,I32096);
  IV  NOT_913(I16168,g3321);
  IV  NOT_914(g26869,g24842);
  IV  NOT_915(g32689,g30825);
  IV  NOT_916(g15824,I17324);
  IV  NOT_917(g20442,g15171);
  IV  NOT_918(g10382,g6958);
  IV  NOT_919(I18912,g15050);
  IV  NOT_920(I22240,g20086);
  IV  NOT_921(g32923,g31021);
  IV  NOT_922(g33451,g32132);
  IV  NOT_923(g19786,g17062);
  IV  NOT_924(I14833,g10142);
  IV  NOT_925(g16659,I17857);
  IV  NOT_926(g12614,g9935);
  IV  NOT_927(g22761,g21024);
  IV  NOT_928(g9280,I13054);
  IV  NOT_929(g10519,g9326);
  IV  NOT_930(g34736,I32904);
  IV  NOT_931(g10176,g44);
  IV  NOT_932(I16479,g10430);
  IV  NOT_933(g27320,I26004);
  IV  NOT_934(g16987,I18135);
  IV  NOT_935(g32688,g30735);
  IV  NOT_936(g32624,g30825);
  IV  NOT_937(I23312,g21681);
  IV  NOT_938(g13279,I15843);
  IV  NOT_939(I16217,g3632);
  IV  NOT_940(I21115,g15714);
  IV  NOT_941(g16658,g14157);
  IV  NOT_942(I22604,g21143);
  IV  NOT_943(g10518,g9311);
  IV  NOT_944(g10154,g2547);
  IV  NOT_945(g12905,g10408);
  IV  NOT_946(g20615,g15509);
  IV  NOT_947(g33246,g32212);
  IV  NOT_948(g9083,g626);
  IV  NOT_949(g23875,g18997);
  IV  NOT_950(g25080,g23742);
  IV  NOT_951(g24116,g21143);
  IV  NOT_952(g14518,I16639);
  IV  NOT_953(g23219,I22316);
  IV  NOT_954(I18051,g13680);
  IV  NOT_955(g30330,I28591);
  IV  NOT_956(g13278,g10738);
  IV  NOT_957(g26709,g25435);
  IV  NOT_958(I29969,g30991);
  IV  NOT_959(g8219,g3731);
  IV  NOT_960(g27565,g26645);
  IV  NOT_961(I17491,g13416);
  IV  NOT_962(I16486,g11204);
  IV  NOT_963(g20041,g15569);
  IV  NOT_964(g9636,g72);
  IV  NOT_965(g22214,g19210);
  IV  NOT_966(g7827,g4688);
  IV  NOT_967(g12122,g9705);
  IV  NOT_968(g20275,g17929);
  IV  NOT_969(g24041,g19968);
  IV  NOT_970(g19998,g15915);
  IV  NOT_971(g8431,g3085);
  IV  NOT_972(g11468,g7624);
  IV  NOT_973(g16644,I17842);
  IV  NOT_974(g13039,I15663);
  IV  NOT_975(g8812,I12805);
  IV  NOT_976(g15426,I17121);
  IV  NOT_977(g22207,I21787);
  IV  NOT_978(g6828,g1300);
  IV  NOT_979(g19672,g16931);
  IV  NOT_980(g34132,g33831);
  IV  NOT_981(g17400,I18333);
  IV  NOT_982(I12890,g4219);
  IV  NOT_983(g29045,g27779);
  IV  NOT_984(g34960,I33218);
  IV  NOT_985(g11038,g8632);
  IV  NOT_986(g16969,g14262);
  IV  NOT_987(g6830,g1389);
  IV  NOT_988(g17013,g14262);
  IV  NOT_989(I18350,g13716);
  IV  NOT_990(g8005,g3025);
  IV  NOT_991(g20237,g17213);
  IV  NOT_992(g21160,g17508);
  IV  NOT_993(g7196,I11860);
  IV  NOT_994(g11815,g7582);
  IV  NOT_995(g8405,I12572);
  IV  NOT_996(g9187,g518);
  IV  NOT_997(g16968,g14238);
  IV  NOT_998(I27552,g28162);
  IV  NOT_999(I15677,g5654);
  IV  NOT_1000(g31859,g29385);
  IV  NOT_1001(I32116,g33937);
  IV  NOT_1002(g20035,g16430);
  IV  NOT_1003(g31825,g29385);
  IV  NOT_1004(g32876,g30735);
  IV  NOT_1005(g32885,g31021);
  IV  NOT_1006(g34161,g33851);
  IV  NOT_1007(g16197,g13861);
  IV  NOT_1008(g24035,g20841);
  IV  NOT_1009(g11677,g7689);
  IV  NOT_1010(g21455,g15426);
  IV  NOT_1011(I12003,g767);
  IV  NOT_1012(g8286,g53);
  IV  NOT_1013(g8765,g3333);
  IV  NOT_1014(g17328,I18313);
  IV  NOT_1015(g31858,g29385);
  IV  NOT_1016(g13975,g11048);
  IV  NOT_1017(g32854,g30735);
  IV  NOT_1018(g7780,g2878);
  IV  NOT_1019(I12779,g4210);
  IV  NOT_1020(g16527,g14048);
  IV  NOT_1021(g25198,g22228);
  IV  NOT_1022(g30259,g28463);
  IV  NOT_1023(g25529,g22763);
  IV  NOT_1024(g14215,g12198);
  IV  NOT_1025(g32511,g30614);
  IV  NOT_1026(g23915,g19277);
  IV  NOT_1027(g32763,g31710);
  IV  NOT_1028(I15937,g11676);
  IV  NOT_1029(I17395,g12952);
  IV  NOT_1030(I28434,g28114);
  IV  NOT_1031(g30087,g29121);
  IV  NOT_1032(g11143,g8032);
  IV  NOT_1033(g19961,g17328);
  IV  NOT_1034(g26810,g25220);
  IV  NOT_1035(I29894,g31771);
  IV  NOT_1036(I14033,g8912);
  IV  NOT_1037(g34471,g34423);
  IV  NOT_1038(g9200,g1548);
  IV  NOT_1039(g25528,g22594);
  IV  NOT_1040(I21934,g21273);
  IV  NOT_1041(g31844,g29385);
  IV  NOT_1042(I31597,g33187);
  IV  NOT_1043(g8733,g3698);
  IV  NOT_1044(g19505,g16349);
  IV  NOT_1045(g23277,I22380);
  IV  NOT_1046(g7018,g5297);
  IV  NOT_1047(g8974,I12930);
  IV  NOT_1048(I11726,g4273);
  IV  NOT_1049(I32237,g34130);
  IV  NOT_1050(I17633,g13258);
  IV  NOT_1051(g32660,g30825);
  IV  NOT_1052(g7418,g2361);
  IV  NOT_1053(I13726,g4537);
  IV  NOT_1054(g9003,g790);
  IV  NOT_1055(g6953,g4157);
  IV  NOT_1056(g7994,I12336);
  IV  NOT_1057(g29997,g29060);
  IV  NOT_1058(g11884,g8125);
  IV  NOT_1059(g21467,g15758);
  IV  NOT_1060(I16676,g10588);
  IV  NOT_1061(g25869,g25250);
  IV  NOT_1062(g10349,g6956);
  IV  NOT_1063(g23494,I22619);
  IV  NOT_1064(g26337,g24818);
  IV  NOT_1065(I32806,g34585);
  IV  NOT_1066(g8796,g4785);
  IV  NOT_1067(I32684,g34430);
  IV  NOT_1068(g32456,g31376);
  IV  NOT_1069(g34244,I32231);
  IV  NOT_1070(I33300,g35001);
  IV  NOT_1071(g20130,g17328);
  IV  NOT_1072(g22683,I22000);
  IV  NOT_1073(g13410,I15921);
  IV  NOT_1074(I12826,g4349);
  IV  NOT_1075(g21037,I20913);
  IV  NOT_1076(g24130,g20998);
  IV  NOT_1077(g32480,g31070);
  IV  NOT_1078(g10083,g2407);
  IV  NOT_1079(g10348,I13762);
  IV  NOT_1080(g32916,g31021);
  IV  NOT_1081(g14348,g10887);
  IV  NOT_1082(g12891,g10399);
  IV  NOT_1083(g8324,g2476);
  IV  NOT_1084(g26792,g25439);
  IV  NOT_1085(g20523,g17821);
  IV  NOT_1086(I16417,g875);
  IV  NOT_1087(I21013,g15806);
  IV  NOT_1088(g32550,g31376);
  IV  NOT_1089(g9637,I13252);
  IV  NOT_1090(g23984,g19210);
  IV  NOT_1091(g18952,g16053);
  IV  NOT_1092(g24165,I23339);
  IV  NOT_1093(g30068,g29157);
  IV  NOT_1094(g34810,I33020);
  IV  NOT_1095(g31227,g29744);
  IV  NOT_1096(g17683,g15027);
  IV  NOT_1097(g23419,g21468);
  IV  NOT_1098(g34068,g33728);
  IV  NOT_1099(g21352,g16322);
  IV  NOT_1100(g13015,g11875);
  IV  NOT_1101(g8540,g3408);
  IV  NOT_1102(g23352,g20924);
  IV  NOT_1103(g25259,I24445);
  IV  NOT_1104(g25225,g23802);
  IV  NOT_1105(g21155,g15656);
  IV  NOT_1106(g34879,I33109);
  IV  NOT_1107(g21418,g17821);
  IV  NOT_1108(g22882,g20391);
  IV  NOT_1109(g28608,g27670);
  IV  NOT_1110(g23418,g21468);
  IV  NOT_1111(g32721,g31021);
  IV  NOT_1112(g20006,g17328);
  IV  NOT_1113(I26466,g26870);
  IV  NOT_1114(I15556,g11928);
  IV  NOT_1115(g32596,g31070);
  IV  NOT_1116(g9223,g1216);
  IV  NOT_1117(g12109,I14967);
  IV  NOT_1118(g19433,g15915);
  IV  NOT_1119(g23170,g20046);
  IV  NOT_1120(g7197,g812);
  IV  NOT_1121(g22407,g19455);
  IV  NOT_1122(g34878,I33106);
  IV  NOT_1123(g19387,g16431);
  IV  NOT_1124(I16762,g5290);
  IV  NOT_1125(g6848,g2417);
  IV  NOT_1126(g7397,g890);
  IV  NOT_1127(I27449,g27737);
  IV  NOT_1128(g15969,I17416);
  IV  NOT_1129(I20846,g16923);
  IV  NOT_1130(g19620,g17296);
  IV  NOT_1131(g12108,I14964);
  IV  NOT_1132(g10139,g136);
  IV  NOT_1133(I15223,g10119);
  IV  NOT_1134(I17612,g13250);
  IV  NOT_1135(I24396,g23453);
  IV  NOT_1136(g6855,g2711);
  IV  NOT_1137(g17414,g14627);
  IV  NOT_1138(g27492,g26598);
  IV  NOT_1139(g8287,g160);
  IV  NOT_1140(I17324,g14119);
  IV  NOT_1141(g9416,g2429);
  IV  NOT_1142(g13223,I15800);
  IV  NOT_1143(g24437,g22654);
  IV  NOT_1144(g25244,g23802);
  IV  NOT_1145(g19343,g16136);
  IV  NOT_1146(g34994,I33282);
  IV  NOT_1147(I17098,g14336);
  IV  NOT_1148(g32773,g31376);
  IV  NOT_1149(g32942,g30825);
  IV  NOT_1150(g9251,I13037);
  IV  NOT_1151(g20703,g15373);
  IV  NOT_1152(g29220,I27576);
  IV  NOT_1153(I11635,g9);
  IV  NOT_1154(g23589,g21468);
  IV  NOT_1155(g10415,g7109);
  IV  NOT_1156(g18422,I19238);
  IV  NOT_1157(g32655,g30614);
  IV  NOT_1158(g8399,g3798);
  IV  NOT_1159(g11110,g8728);
  IV  NOT_1160(g29911,g28780);
  IV  NOT_1161(g19369,g15995);
  IV  NOT_1162(g33377,I30901);
  IV  NOT_1163(g34425,I32446);
  IV  NOT_1164(g12381,I15223);
  IV  NOT_1165(g23524,g21562);
  IV  NOT_1166(g27091,g26725);
  IV  NOT_1167(g28184,I26705);
  IV  NOT_1168(g32670,g30673);
  IV  NOT_1169(g33120,I30686);
  IV  NOT_1170(I12026,g344);
  IV  NOT_1171(I21100,g16284);
  IV  NOT_1172(g8898,g676);
  IV  NOT_1173(g20600,g15348);
  IV  NOT_1174(I16117,g10430);
  IV  NOT_1175(g34919,I33149);
  IV  NOT_1176(g19368,g16326);
  IV  NOT_1177(I32222,g34118);
  IV  NOT_1178(g20781,I20840);
  IV  NOT_1179(g16877,I18071);
  IV  NOT_1180(g23477,g21468);
  IV  NOT_1181(g32734,g31710);
  IV  NOT_1182(g33645,I31477);
  IV  NOT_1183(g22759,g19857);
  IV  NOT_1184(I17140,g13835);
  IV  NOT_1185(g26817,g25242);
  IV  NOT_1186(g7631,g74);
  IV  NOT_1187(g34918,I33146);
  IV  NOT_1188(g17584,g14773);
  IV  NOT_1189(I26693,g27930);
  IV  NOT_1190(g10664,g8928);
  IV  NOT_1191(I20929,g17663);
  IV  NOT_1192(g32839,g30735);
  IV  NOT_1193(g32930,g31021);
  IV  NOT_1194(g20372,g17847);
  IV  NOT_1195(g30079,g29097);
  IV  NOT_1196(g19412,g16489);
  IV  NOT_1197(g7257,I11903);
  IV  NOT_1198(g22758,g20330);
  IV  NOT_1199(g24372,g22885);
  IV  NOT_1200(g16695,g14454);
  IV  NOT_1201(g25171,g22228);
  IV  NOT_1202(g20175,I20433);
  IV  NOT_1203(g7301,g925);
  IV  NOT_1204(I16747,g12729);
  IV  NOT_1205(g8291,I12503);
  IV  NOT_1206(g11373,g7566);
  IV  NOT_1207(g23864,g19210);
  IV  NOT_1208(g25886,g24537);
  IV  NOT_1209(g23022,g20283);
  IV  NOT_1210(g32667,g30825);
  IV  NOT_1211(g32694,g31376);
  IV  NOT_1212(g32838,g31376);
  IV  NOT_1213(I31550,g33204);
  IV  NOT_1214(g33698,I31539);
  IV  NOT_1215(g24175,I23369);
  IV  NOT_1216(g29147,I27449);
  IV  NOT_1217(g32965,g31710);
  IV  NOT_1218(g12840,g10356);
  IV  NOT_1219(g6818,g976);
  IV  NOT_1220(g17759,g14864);
  IV  NOT_1221(g6867,I11685);
  IV  NOT_1222(g16526,g13898);
  IV  NOT_1223(g23749,g18997);
  IV  NOT_1224(I15800,g11607);
  IV  NOT_1225(g15714,I17228);
  IV  NOT_1226(g9880,g5787);
  IV  NOT_1227(g23313,g21070);
  IV  NOT_1228(g25994,g24575);
  IV  NOT_1229(g8344,I12523);
  IV  NOT_1230(g9537,g1748);
  IV  NOT_1231(g29950,g28896);
  IV  NOT_1232(g24063,g20014);
  IV  NOT_1233(g17758,g14861);
  IV  NOT_1234(g26656,g25495);
  IV  NOT_1235(g20516,I20609);
  IV  NOT_1236(g10554,g8974);
  IV  NOT_1237(g18905,g16077);
  IV  NOT_1238(g24137,g20998);
  IV  NOT_1239(g32487,g30825);
  IV  NOT_1240(g24516,g22670);
  IV  NOT_1241(g7751,g1521);
  IV  NOT_1242(g23285,g20887);
  IV  NOT_1243(g26680,g25300);
  IV  NOT_1244(g32619,g30614);
  IV  NOT_1245(g8259,g2217);
  IV  NOT_1246(g21305,g15758);
  IV  NOT_1247(g21053,g15373);
  IV  NOT_1248(g32502,g31070);
  IV  NOT_1249(g14609,I16724);
  IV  NOT_1250(g15979,I17420);
  IV  NOT_1251(g10200,g2138);
  IV  NOT_1252(g23305,g20391);
  IV  NOT_1253(g32557,g31376);
  IV  NOT_1254(g13334,g11048);
  IV  NOT_1255(g29151,g27858);
  IV  NOT_1256(g29172,g27020);
  IV  NOT_1257(I24787,g24266);
  IV  NOT_1258(g9978,g2756);
  IV  NOT_1259(g30322,g28431);
  IV  NOT_1260(g10608,g9155);
  IV  NOT_1261(g29996,g28962);
  IV  NOT_1262(I12811,g4340);
  IV  NOT_1263(g10115,g2283);
  IV  NOT_1264(I16639,g4000);
  IV  NOT_1265(g21466,g15509);
  IV  NOT_1266(g32618,g31154);
  IV  NOT_1267(I18662,g6322);
  IV  NOT_1268(g8088,g1554);
  IV  NOT_1269(g6975,g4507);
  IV  NOT_1270(g9417,I13124);
  IV  NOT_1271(g34159,I32116);
  IV  NOT_1272(g11762,g7964);
  IV  NOT_1273(g7041,g5644);
  IV  NOT_1274(g9935,I13483);
  IV  NOT_1275(I13606,g74);
  IV  NOT_1276(g11964,g9154);
  IV  NOT_1277(g21036,I20910);
  IV  NOT_1278(g7441,g862);
  IV  NOT_1279(g20209,g17821);
  IV  NOT_1280(g33661,I31497);
  IV  NOT_1281(g33895,I31751);
  IV  NOT_1282(g9982,g3976);
  IV  NOT_1283(g21177,I20957);
  IV  NOT_1284(g21560,g17873);
  IV  NOT_1285(g16077,I17456);
  IV  NOT_1286(g9234,g5170);
  IV  NOT_1287(I15587,g11985);
  IV  NOT_1288(g32469,g30673);
  IV  NOT_1289(I27368,g27881);
  IV  NOT_1290(I18482,g13350);
  IV  NOT_1291(g20208,g17533);
  IV  NOT_1292(g14745,g12423);
  IV  NOT_1293(g13216,g10939);
  IV  NOT_1294(g17141,I18191);
  IV  NOT_1295(I11750,g4474);
  IV  NOT_1296(I18248,g12938);
  IV  NOT_1297(g19379,g17327);
  IV  NOT_1298(g26631,g25467);
  IV  NOT_1299(g12862,g10370);
  IV  NOT_1300(g17652,g15033);
  IV  NOT_1301(g34656,I32770);
  IV  NOT_1302(g8215,I12451);
  IV  NOT_1303(g30295,I28540);
  IV  NOT_1304(g22332,I21838);
  IV  NOT_1305(g9542,g2173);
  IV  NOT_1306(I16391,g859);
  IV  NOT_1307(g26364,I25327);
  IV  NOT_1308(g32468,g30614);
  IV  NOT_1309(g6821,I11655);
  IV  NOT_1310(I18003,g13638);
  IV  NOT_1311(g19050,I19759);
  IV  NOT_1312(g34680,I32820);
  IV  NOT_1313(g8951,g554);
  IV  NOT_1314(g16689,g13923);
  IV  NOT_1315(g34144,I32093);
  IV  NOT_1316(g34823,I33037);
  IV  NOT_1317(g20542,g17873);
  IV  NOT_1318(g16923,I18089);
  IV  NOT_1319(g20453,I20584);
  IV  NOT_1320(g16280,g13330);
  IV  NOT_1321(g6984,g4709);
  IV  NOT_1322(g32038,g30934);
  IV  NOT_1323(g24021,g20841);
  IV  NOT_1324(g28241,g27064);
  IV  NOT_1325(g29318,g29029);
  IV  NOT_1326(g16688,g14045);
  IV  NOT_1327(g16624,I17814);
  IV  NOT_1328(g22406,g19506);
  IV  NOT_1329(g8114,g3522);
  IV  NOT_1330(g10184,g4486);
  IV  NOT_1331(g12040,I14902);
  IV  NOT_1332(I16579,g10981);
  IV  NOT_1333(g16300,I17626);
  IV  NOT_1334(g19386,g16431);
  IV  NOT_1335(g10805,I14046);
  IV  NOT_1336(I22785,g18940);
  IV  NOT_1337(g20913,g15373);
  IV  NOT_1338(I18778,g6704);
  IV  NOT_1339(g34336,g34112);
  IV  NOT_1340(g32815,g30937);
  IV  NOT_1341(g14184,g12381);
  IV  NOT_1342(g19603,g16349);
  IV  NOT_1343(g19742,g17096);
  IV  NOT_1344(g13117,g10981);
  IV  NOT_1345(g17135,g14297);
  IV  NOT_1346(g12904,g10410);
  IV  NOT_1347(g20614,g15426);
  IV  NOT_1348(g32601,g31376);
  IV  NOT_1349(I15569,g11965);
  IV  NOT_1350(g9554,g5105);
  IV  NOT_1351(g20436,I20569);
  IV  NOT_1352(g23874,g18997);
  IV  NOT_1353(g8870,I12837);
  IV  NOT_1354(g32677,g30673);
  IV  NOT_1355(g33127,g31950);
  IV  NOT_1356(g25322,I24497);
  IV  NOT_1357(I31694,g33176);
  IV  NOT_1358(I32834,g34472);
  IV  NOT_1359(g32975,I30537);
  IV  NOT_1360(g21693,I21254);
  IV  NOT_1361(g20607,g17955);
  IV  NOT_1362(g13569,g10951);
  IV  NOT_1363(g8650,g4664);
  IV  NOT_1364(I12896,g4229);
  IV  NOT_1365(g20320,g17015);
  IV  NOT_1366(I18647,g5320);
  IV  NOT_1367(g20073,g16540);
  IV  NOT_1368(I28832,g30301);
  IV  NOT_1369(I33131,g34906);
  IV  NOT_1370(g30017,g29085);
  IV  NOT_1371(g20274,g17847);
  IV  NOT_1372(g9213,I13020);
  IV  NOT_1373(g24073,g21127);
  IV  NOT_1374(g20530,g15509);
  IV  NOT_1375(g21665,I21226);
  IV  NOT_1376(g25158,g22228);
  IV  NOT_1377(I21744,g19338);
  IV  NOT_1378(g20593,g15277);
  IV  NOT_1379(I17754,g13494);
  IV  NOT_1380(g23665,g21562);
  IV  NOT_1381(g25783,g25250);
  IV  NOT_1382(I17355,g14591);
  IV  NOT_1383(g32937,g31021);
  IV  NOT_1384(g19429,g16489);
  IV  NOT_1385(I23345,g23320);
  IV  NOT_1386(g33385,g32038);
  IV  NOT_1387(I21849,g19620);
  IV  NOT_1388(g29044,g27742);
  IV  NOT_1389(g10761,g8411);
  IV  NOT_1390(g7411,g2040);
  IV  NOT_1391(g25561,g22550);
  IV  NOT_1392(g18891,g16053);
  IV  NOT_1393(g20565,g18008);
  IV  NOT_1394(I31619,g33212);
  IV  NOT_1395(I15814,g11129);
  IV  NOT_1396(g24122,g20857);
  IV  NOT_1397(I23399,g23450);
  IV  NOT_1398(g8136,g269);
  IV  NOT_1399(g19730,g17062);
  IV  NOT_1400(g19428,g16090);
  IV  NOT_1401(g12183,I15033);
  IV  NOT_1402(g9902,g100);
  IV  NOT_1403(I18233,g14639);
  IV  NOT_1404(g33354,g32329);
  IV  NOT_1405(I33210,g34943);
  IV  NOT_1406(g32791,g31672);
  IV  NOT_1407(g23476,g21468);
  IV  NOT_1408(g23485,g20785);
  IV  NOT_1409(I25555,g25241);
  IV  NOT_1410(g31824,g29385);
  IV  NOT_1411(g32884,g30825);
  IV  NOT_1412(g33888,g33346);
  IV  NOT_1413(g8594,g3849);
  IV  NOT_1414(g19765,g16897);
  IV  NOT_1415(g6756,I11623);
  IV  NOT_1416(g24034,g19968);
  IV  NOT_1417(g7074,I11801);
  IV  NOT_1418(g11772,I14623);
  IV  NOT_1419(g10400,g7002);
  IV  NOT_1420(g20641,g15509);
  IV  NOT_1421(g26816,g25260);
  IV  NOT_1422(g21454,g15373);
  IV  NOT_1423(I33279,g34986);
  IV  NOT_1424(g23555,I22692);
  IV  NOT_1425(I32607,g34358);
  IV  NOT_1426(g7474,I11980);
  IV  NOT_1427(g17221,I18245);
  IV  NOT_1428(g19690,g16826);
  IV  NOT_1429(g30309,g28959);
  IV  NOT_1430(g7992,g5008);
  IV  NOT_1431(g9490,g2563);
  IV  NOT_1432(I14563,g802);
  IV  NOT_1433(g16511,g14130);
  IV  NOT_1434(g9166,g837);
  IV  NOT_1435(g20153,g16782);
  IV  NOT_1436(g23570,g18833);
  IV  NOT_1437(I32274,g34195);
  IV  NOT_1438(g23914,g19210);
  IV  NOT_1439(g32479,g30735);
  IV  NOT_1440(g32666,g31376);
  IV  NOT_1441(I13483,g6035);
  IV  NOT_1442(g11293,g7527);
  IV  NOT_1443(g24153,I23303);
  IV  NOT_1444(I31469,g33388);
  IV  NOT_1445(g6904,g3494);
  IV  NOT_1446(g32363,I29891);
  IV  NOT_1447(I12112,g794);
  IV  NOT_1448(g12872,g10379);
  IV  NOT_1449(g13638,I16057);
  IV  NOT_1450(g34308,g34088);
  IV  NOT_1451(g9056,g3017);
  IV  NOT_1452(g23907,g19074);
  IV  NOT_1453(g32478,g31376);
  IV  NOT_1454(g32015,I29571);
  IV  NOT_1455(g19504,g16349);
  IV  NOT_1456(g9456,g6073);
  IV  NOT_1457(g33931,I31807);
  IV  NOT_1458(I32464,g34245);
  IV  NOT_1459(g8228,g3835);
  IV  NOT_1460(g9529,g6561);
  IV  NOT_1461(g7863,g1249);
  IV  NOT_1462(g20136,I20399);
  IV  NOT_1463(g20635,g18008);
  IV  NOT_1464(I27742,g28819);
  IV  NOT_1465(g13416,I15929);
  IV  NOT_1466(g25017,g23699);
  IV  NOT_1467(I25567,g25272);
  IV  NOT_1468(I25594,g25531);
  IV  NOT_1469(I18897,g16738);
  IV  NOT_1470(g24136,g20857);
  IV  NOT_1471(g32486,g30735);
  IV  NOT_1472(I13326,g66);
  IV  NOT_1473(g23239,g21308);
  IV  NOT_1474(g33426,g32017);
  IV  NOT_1475(g11841,g9800);
  IV  NOT_1476(g9155,I12997);
  IV  NOT_1477(I14395,g3654);
  IV  NOT_1478(g6841,g2145);
  IV  NOT_1479(I17420,g13394);
  IV  NOT_1480(g23567,g21562);
  IV  NOT_1481(g32556,g31554);
  IV  NOT_1482(I32797,g34581);
  IV  NOT_1483(I14899,g10198);
  IV  NOT_1484(g8033,g157);
  IV  NOT_1485(g23238,g20924);
  IV  NOT_1486(g11510,g7633);
  IV  NOT_1487(g13510,I15981);
  IV  NOT_1488(g17812,I18810);
  IV  NOT_1489(g34816,I33030);
  IV  NOT_1490(I20647,g17010);
  IV  NOT_1491(g32580,g30825);
  IV  NOT_1492(g9698,g2181);
  IV  NOT_1493(g28441,g27629);
  IV  NOT_1494(g26260,g24759);
  IV  NOT_1495(I14633,g9340);
  IV  NOT_1496(g9964,g126);
  IV  NOT_1497(I13252,g6751);
  IV  NOT_1498(g20164,g16826);
  IV  NOT_1499(g34985,I33255);
  IV  NOT_1500(I20999,g16709);
  IV  NOT_1501(g23941,g19074);
  IV  NOT_1502(g18091,I18879);
  IV  NOT_1503(g19128,I19778);
  IV  NOT_1504(g23382,g20682);
  IV  NOT_1505(g24164,I23336);
  IV  NOT_1506(g25289,g22228);
  IV  NOT_1507(g21176,I20954);
  IV  NOT_1508(g21185,g15277);
  IV  NOT_1509(g23519,g21468);
  IV  NOT_1510(I27730,g28752);
  IV  NOT_1511(g12047,g9591);
  IV  NOT_1512(g16307,I17633);
  IV  NOT_1513(g13835,I16150);
  IV  NOT_1514(g34954,I33210);
  IV  NOT_1515(g13014,g11872);
  IV  NOT_1516(g25023,g22457);
  IV  NOT_1517(g24891,g23231);
  IV  NOT_1518(I33143,g34903);
  IV  NOT_1519(g19626,g17409);
  IV  NOT_1520(g25288,g22228);
  IV  NOT_1521(g25224,g22763);
  IV  NOT_1522(I20233,g17487);
  IV  NOT_1523(g16721,g14072);
  IV  NOT_1524(I12793,g4578);
  IV  NOT_1525(g23518,g21070);
  IV  NOT_1526(g23154,I22264);
  IV  NOT_1527(g26488,I25366);
  IV  NOT_1528(g26424,I25356);
  IV  NOT_1529(g20575,g17929);
  IV  NOT_1530(g31860,I29438);
  IV  NOT_1531(g13007,g11852);
  IV  NOT_1532(g25308,g22763);
  IV  NOT_1533(g8195,g1783);
  IV  NOT_1534(g8137,g411);
  IV  NOT_1535(g32922,g31710);
  IV  NOT_1536(g8891,g582);
  IV  NOT_1537(g19533,g16261);
  IV  NOT_1538(g24474,g23620);
  IV  NOT_1539(g20711,g15509);
  IV  NOT_1540(I16193,g3281);
  IV  NOT_1541(g16431,I17675);
  IV  NOT_1542(I27549,g28161);
  IV  NOT_1543(g27051,I25779);
  IV  NOT_1544(g32531,g31070);
  IV  NOT_1545(I13847,g7266);
  IV  NOT_1546(I31791,g33354);
  IV  NOT_1547(g20327,g15224);
  IV  NOT_1548(g23935,g19210);
  IV  NOT_1549(g24711,g23139);
  IV  NOT_1550(g34669,I32791);
  IV  NOT_1551(g26830,g24411);
  IV  NOT_1552(g27592,g26715);
  IV  NOT_1553(g12051,g9595);
  IV  NOT_1554(g20537,g15345);
  IV  NOT_1555(g24109,g21143);
  IV  NOT_1556(g32740,g31672);
  IV  NOT_1557(g15885,I17374);
  IV  NOT_1558(g8807,g79);
  IV  NOT_1559(g11615,g6875);
  IV  NOT_1560(g9619,g5845);
  IV  NOT_1561(g17507,g15030);
  IV  NOT_1562(I24331,g22976);
  IV  NOT_1563(g34668,I32788);
  IV  NOT_1564(g13116,g10935);
  IV  NOT_1565(g16773,g14021);
  IV  NOT_1566(I18148,g13526);
  IV  NOT_1567(g24108,g20998);
  IV  NOT_1568(I28162,g28803);
  IV  NOT_1569(g32186,I29720);
  IV  NOT_1570(g34392,g34202);
  IV  NOT_1571(g32676,g30614);
  IV  NOT_1572(g32685,g31528);
  IV  NOT_1573(g33659,I31491);
  IV  NOT_1574(g28399,g27074);
  IV  NOT_1575(g30195,I28434);
  IV  NOT_1576(g7400,g911);
  IV  NOT_1577(g8859,g772);
  IV  NOT_1578(g32953,g31327);
  IV  NOT_1579(g19737,g17015);
  IV  NOT_1580(g11720,I14589);
  IV  NOT_1581(g20283,I20529);
  IV  NOT_1582(g6811,g714);
  IV  NOT_1583(g34195,I32150);
  IV  NOT_1584(g20606,g17955);
  IV  NOT_1585(g33250,g32186);
  IV  NOT_1586(g16655,g14151);
  IV  NOT_1587(g10882,g7601);
  IV  NOT_1588(I18104,g13177);
  IV  NOT_1589(g10414,g7092);
  IV  NOT_1590(I13634,g79);
  IV  NOT_1591(g31658,I29242);
  IV  NOT_1592(I13872,g7474);
  IV  NOT_1593(g13041,I15667);
  IV  NOT_1594(g32654,g31070);
  IV  NOT_1595(g9843,g4311);
  IV  NOT_1596(g33658,g33080);
  IV  NOT_1597(g16180,g13437);
  IV  NOT_1598(g30016,g29049);
  IV  NOT_1599(g9989,g5077);
  IV  NOT_1600(I24448,g22923);
  IV  NOT_1601(g11430,g7617);
  IV  NOT_1602(g22541,I21911);
  IV  NOT_1603(g34559,g34384);
  IV  NOT_1604(g12350,I15190);
  IV  NOT_1605(g10407,g7063);
  IV  NOT_1606(g32800,g31021);
  IV  NOT_1607(g32936,g31710);
  IV  NOT_1608(g19697,g16886);
  IV  NOT_1609(I31486,g33197);
  IV  NOT_1610(g23215,g20785);
  IV  NOT_1611(g12820,g10233);
  IV  NOT_1612(I17699,g13416);
  IV  NOT_1613(g23501,g20924);
  IV  NOT_1614(g6874,g3143);
  IV  NOT_1615(I29965,g31189);
  IV  NOT_1616(I32109,g33631);
  IV  NOT_1617(I21033,g17221);
  IV  NOT_1618(g20381,g17955);
  IV  NOT_1619(g8342,I12519);
  IV  NOT_1620(g11237,I14305);
  IV  NOT_1621(g9834,g2579);
  IV  NOT_1622(g9971,g2093);
  IV  NOT_1623(I21234,g16540);
  IV  NOT_1624(g24982,g22763);
  IV  NOT_1625(g26679,g25385);
  IV  NOT_1626(g34830,I33044);
  IV  NOT_1627(g34893,I33119);
  IV  NOT_1628(g9686,g73);
  IV  NOT_1629(g22359,g19495);
  IV  NOT_1630(g8255,g2028);
  IV  NOT_1631(g17473,g14841);
  IV  NOT_1632(g20091,g17328);
  IV  NOT_1633(I22366,g19757);
  IV  NOT_1634(g24091,g20720);
  IV  NOT_1635(g7183,g4608);
  IV  NOT_1636(g8481,I12618);
  IV  NOT_1637(I12128,g4253);
  IV  NOT_1638(g17789,g14321);
  IV  NOT_1639(g29956,I28185);
  IV  NOT_1640(g29385,g28180);
  IV  NOT_1641(g34544,I32613);
  IV  NOT_1642(g15480,I17125);
  IV  NOT_1643(I26664,g27708);
  IV  NOT_1644(g22358,g19801);
  IV  NOT_1645(g32762,g31672);
  IV  NOT_1646(g9598,g2571);
  IV  NOT_1647(g24174,I23366);
  IV  NOT_1648(g8097,g3029);
  IV  NOT_1649(g25260,I24448);
  IV  NOT_1650(g32964,g31672);
  IV  NOT_1651(g29980,g28935);
  IV  NOT_1652(g7779,g1413);
  IV  NOT_1653(g34713,I32871);
  IV  NOT_1654(g8497,g3436);
  IV  NOT_1655(g13142,g10632);
  IV  NOT_1656(g21349,g15758);
  IV  NOT_1657(g8154,g3139);
  IV  NOT_1658(I28591,g29371);
  IV  NOT_1659(g17325,I18304);
  IV  NOT_1660(g8354,g4815);
  IV  NOT_1661(g18948,g15800);
  IV  NOT_1662(g7023,g5445);
  IV  NOT_1663(g31855,g29385);
  IV  NOT_1664(g10206,g4489);
  IV  NOT_1665(g14441,I16590);
  IV  NOT_1666(g14584,g11048);
  IV  NOT_1667(g9321,g5863);
  IV  NOT_1668(g7423,g2433);
  IV  NOT_1669(g9670,g5022);
  IV  NOT_1670(I22547,g20720);
  IV  NOT_1671(g25195,g22763);
  IV  NOT_1672(g16487,I17695);
  IV  NOT_1673(g23906,g19074);
  IV  NOT_1674(g26093,g24814);
  IV  NOT_1675(g30610,I28872);
  IV  NOT_1676(g18904,g16053);
  IV  NOT_1677(g32587,g30735);
  IV  NOT_1678(g15085,I17008);
  IV  NOT_1679(I32982,g34749);
  IV  NOT_1680(g23284,g20785);
  IV  NOT_1681(g19445,g15915);
  IV  NOT_1682(g10725,g7846);
  IV  NOT_1683(g21304,g17367);
  IV  NOT_1684(g25525,g22550);
  IV  NOT_1685(g34042,g33674);
  IV  NOT_1686(g25424,g23800);
  IV  NOT_1687(I20433,g16234);
  IV  NOT_1688(g23304,g20785);
  IV  NOT_1689(g25016,g23666);
  IV  NOT_1690(g6978,g4616);
  IV  NOT_1691(I33179,g34893);
  IV  NOT_1692(g7161,I11843);
  IV  NOT_1693(g19499,g16782);
  IV  NOT_1694(g17121,g14321);
  IV  NOT_1695(g7361,g1874);
  IV  NOT_1696(g22682,g19379);
  IV  NOT_1697(g10114,g2116);
  IV  NOT_1698(g20192,g17268);
  IV  NOT_1699(g9253,g5037);
  IV  NOT_1700(I16821,g5983);
  IV  NOT_1701(I17661,g13329);
  IV  NOT_1702(g27929,I26448);
  IV  NOT_1703(g25558,g22594);
  IV  NOT_1704(g23566,g21562);
  IV  NOT_1705(g32909,g30614);
  IV  NOT_1706(g10082,g2375);
  IV  NOT_1707(g32543,g31376);
  IV  NOT_1708(g34270,g34159);
  IV  NOT_1709(I27232,g27993);
  IV  NOT_1710(g19498,g16752);
  IV  NOT_1711(g34188,g33875);
  IV  NOT_1712(g7051,I11793);
  IV  NOT_1713(g10107,I13606);
  IV  NOT_1714(g22173,I21757);
  IV  NOT_1715(g34124,g33819);
  IV  NOT_1716(g9909,g1978);
  IV  NOT_1717(g12929,g12550);
  IV  NOT_1718(g25830,g24485);
  IV  NOT_1719(g27583,g26686);
  IV  NOT_1720(g20663,g15373);
  IV  NOT_1721(g27928,g26810);
  IV  NOT_1722(g25893,g24541);
  IV  NOT_1723(g8783,I12761);
  IV  NOT_1724(g7451,g2070);
  IV  NOT_1725(g32908,g31327);
  IV  NOT_1726(g6982,g4531);
  IV  NOT_1727(g7327,g2165);
  IV  NOT_1728(g24522,g22689);
  IV  NOT_1729(g33894,I31748);
  IV  NOT_1730(g11165,I14222);
  IV  NOT_1731(g8112,g3419);
  IV  NOT_1732(g8218,g3490);
  IV  NOT_1733(g34939,g34922);
  IV  NOT_1734(g9740,g5821);
  IV  NOT_1735(g8267,g2342);
  IV  NOT_1736(g25544,g22594);
  IV  NOT_1737(g32569,g30673);
  IV  NOT_1738(g34383,I32388);
  IV  NOT_1739(g29190,g27046);
  IV  NOT_1740(I32840,g34480);
  IV  NOT_1741(g17291,I18276);
  IV  NOT_1742(g14744,g12578);
  IV  NOT_1743(g16286,I17615);
  IV  NOT_1744(g21139,g15634);
  IV  NOT_1745(g21653,g17663);
  IV  NOT_1746(g26837,g24869);
  IV  NOT_1747(g7633,I12120);
  IV  NOT_1748(g34938,g34920);
  IV  NOT_1749(g23653,I22788);
  IV  NOT_1750(g9552,g3654);
  IV  NOT_1751(g15655,g13202);
  IV  NOT_1752(I31800,g33164);
  IV  NOT_1753(g10399,g7017);
  IV  NOT_1754(g32568,g31170);
  IV  NOT_1755(g32747,g30825);
  IV  NOT_1756(I18310,g12978);
  IV  NOT_1757(I20369,g17690);
  IV  NOT_1758(g18062,I18872);
  IV  NOT_1759(g21138,g15634);
  IV  NOT_1760(g24483,I23688);
  IV  NOT_1761(g19432,g15885);
  IV  NOT_1762(I19837,g1399);
  IV  NOT_1763(g30065,g29049);
  IV  NOT_1764(I11820,g3869);
  IV  NOT_1765(g23138,g20453);
  IV  NOT_1766(I26799,g27660);
  IV  NOT_1767(g20553,g17929);
  IV  NOT_1768(g31819,g29385);
  IV  NOT_1769(g8676,g4821);
  IV  NOT_1770(I15727,g10981);
  IV  NOT_1771(I32192,g33628);
  IV  NOT_1772(g10398,g6999);
  IV  NOT_1773(I18379,g13012);
  IV  NOT_1774(g14398,I16555);
  IV  NOT_1775(g10141,I13634);
  IV  NOT_1776(g29211,I27549);
  IV  NOT_1777(g10652,g7601);
  IV  NOT_1778(g10804,g9772);
  IV  NOT_1779(g6800,g203);
  IV  NOT_1780(I13152,g6746);
  IV  NOT_1781(g9687,I13287);
  IV  NOT_1782(g31818,g29385);
  IV  NOT_1783(g32814,g31021);
  IV  NOT_1784(g20326,g18008);
  IV  NOT_1785(g23333,g20785);
  IV  NOT_1786(g13222,g10590);
  IV  NOT_1787(g19753,g16987);
  IV  NOT_1788(g16601,I17783);
  IV  NOT_1789(g17760,I18752);
  IV  NOT_1790(g16677,I17879);
  IV  NOT_1791(I22889,g18926);
  IV  NOT_1792(g20536,g18065);
  IV  NOT_1793(g20040,g17271);
  IV  NOT_1794(g13437,I15937);
  IV  NOT_1795(I20412,g16213);
  IV  NOT_1796(g32751,g31327);
  IV  NOT_1797(g32807,g31021);
  IV  NOT_1798(g32772,g31327);
  IV  NOT_1799(g28463,I26952);
  IV  NOT_1800(g32974,g30937);
  IV  NOT_1801(g8830,g767);
  IV  NOT_1802(g24040,g19919);
  IV  NOT_1803(g7753,I12183);
  IV  NOT_1804(g20702,g17955);
  IV  NOT_1805(g30218,g28918);
  IV  NOT_1806(g25188,g23909);
  IV  NOT_1807(g32639,g31070);
  IV  NOT_1808(g20904,g17433);
  IV  NOT_1809(I17956,g14562);
  IV  NOT_1810(g23963,g19147);
  IV  NOT_1811(g19650,g16971);
  IV  NOT_1812(g28033,g26365);
  IV  NOT_1813(g8592,g3805);
  IV  NOT_1814(g7072,g6199);
  IV  NOT_1815(g14332,I16492);
  IV  NOT_1816(I11691,g36);
  IV  NOT_1817(I28540,g28954);
  IV  NOT_1818(g32638,g30825);
  IV  NOT_1819(g7472,g6329);
  IV  NOT_1820(g19529,g16349);
  IV  NOT_1821(g12640,I15382);
  IV  NOT_1822(I15600,g10430);
  IV  NOT_1823(g22927,I22128);
  IV  NOT_1824(g9860,g5417);
  IV  NOT_1825(g10406,g7046);
  IV  NOT_1826(I24228,g22409);
  IV  NOT_1827(g20564,g15373);
  IV  NOT_1828(g10361,g6841);
  IV  NOT_1829(I25576,g25296);
  IV  NOT_1830(g7443,g914);
  IV  NOT_1831(g8703,I12709);
  IV  NOT_1832(g14406,g12249);
  IV  NOT_1833(g19528,g16349);
  IV  NOT_1834(g19696,g17015);
  IV  NOT_1835(g34160,I32119);
  IV  NOT_1836(g25267,g22228);
  IV  NOT_1837(g19330,g17326);
  IV  NOT_1838(I17181,g13745);
  IV  NOT_1839(I17671,g13280);
  IV  NOT_1840(I29363,g30218);
  IV  NOT_1841(g23585,g21070);
  IV  NOT_1842(g32841,g31672);
  IV  NOT_1843(g11236,g8357);
  IV  NOT_1844(I21291,g18273);
  IV  NOT_1845(g7116,g22);
  IV  NOT_1846(g22649,g19063);
  IV  NOT_1847(g10500,I13875);
  IV  NOT_1848(g27881,I26430);
  IV  NOT_1849(g19365,g16249);
  IV  NOT_1850(g20673,g15277);
  IV  NOT_1851(g32510,g31194);
  IV  NOT_1852(g9691,g1706);
  IV  NOT_1853(g31801,g29385);
  IV  NOT_1854(I15821,g11143);
  IV  NOT_1855(I12056,g2748);
  IV  NOT_1856(g24183,I23393);
  IV  NOT_1857(I32904,g34708);
  IV  NOT_1858(g14833,g11405);
  IV  NOT_1859(g19869,g16540);
  IV  NOT_1860(g21609,g18008);
  IV  NOT_1861(g19960,g17433);
  IV  NOT_1862(g23609,g21611);
  IV  NOT_1863(g24397,g22908);
  IV  NOT_1864(g29339,g28274);
  IV  NOT_1865(g12881,g10388);
  IV  NOT_1866(g7565,I12046);
  IV  NOT_1867(g22903,g20330);
  IV  NOT_1868(g13175,g10909);
  IV  NOT_1869(g34915,I33137);
  IV  NOT_1870(I16593,g10498);
  IV  NOT_1871(I25115,g25322);
  IV  NOT_1872(g32579,g30735);
  IV  NOT_1873(g8068,g3457);
  IV  NOT_1874(I13020,g6750);
  IV  NOT_1875(I32621,g34335);
  IV  NOT_1876(g23312,g21070);
  IV  NOT_1877(I31569,g33197);
  IV  NOT_1878(I28301,g29042);
  IV  NOT_1879(g25219,I24393);
  IV  NOT_1880(I27271,g27998);
  IV  NOT_1881(g21608,g17955);
  IV  NOT_1882(g24062,g19968);
  IV  NOT_1883(g17649,I18614);
  IV  NOT_1884(g20509,g15277);
  IV  NOT_1885(g23608,g21611);
  IV  NOT_1886(g34201,I32158);
  IV  NOT_1887(g9607,g5046);
  IV  NOT_1888(g24509,g22689);
  IV  NOT_1889(g32578,g31376);
  IV  NOT_1890(g32835,g31710);
  IV  NOT_1891(g33695,g33187);
  IV  NOT_1892(g34277,I32274);
  IV  NOT_1893(g25218,g23949);
  IV  NOT_1894(g9962,g6519);
  IV  NOT_1895(g11790,I14630);
  IV  NOT_1896(g14004,g11149);
  IV  NOT_1897(g17648,g15024);
  IV  NOT_1898(g20508,g15277);
  IV  NOT_1899(g9158,g513);
  IV  NOT_1900(g27662,I26296);
  IV  NOT_1901(g17491,g12983);
  IV  NOT_1902(g22981,g20283);
  IV  NOT_1903(g20634,g15373);
  IV  NOT_1904(I21029,g15816);
  IV  NOT_1905(g21052,g15373);
  IV  NOT_1906(g28163,I26682);
  IV  NOT_1907(g8677,g4854);
  IV  NOT_1908(g25837,g25064);
  IV  NOT_1909(g7533,g1306);
  IV  NOT_1910(g19709,g16987);
  IV  NOT_1911(g32586,g31376);
  IV  NOT_1912(I22211,g21463);
  IV  NOT_1913(g9506,g5774);
  IV  NOT_1914(g17604,I18555);
  IV  NOT_1915(g34595,I32693);
  IV  NOT_1916(g7697,g4087);
  IV  NOT_1917(g10613,g10233);
  IV  NOT_1918(g23745,g20900);
  IV  NOT_1919(I18504,g5283);
  IV  NOT_1920(I22024,g19350);
  IV  NOT_1921(g32442,g31213);
  IV  NOT_1922(I31814,g33149);
  IV  NOT_1923(g19471,g16449);
  IV  NOT_1924(g30037,g29121);
  IV  NOT_1925(g12890,g10397);
  IV  NOT_1926(g16580,I17754);
  IV  NOT_1927(g23813,g18997);
  IV  NOT_1928(g7596,I12070);
  IV  NOT_1929(I31751,g33228);
  IV  NOT_1930(I31807,g33149);
  IV  NOT_1931(g16223,g13437);
  IV  NOT_1932(g10273,I13708);
  IV  NOT_1933(g33457,I30989);
  IV  NOT_1934(I32062,g33653);
  IV  NOT_1935(I12199,g6215);
  IV  NOT_1936(g10106,g16);
  IV  NOT_1937(g9311,g5523);
  IV  NOT_1938(I11743,g4564);
  IV  NOT_1939(g22845,g20682);
  IV  NOT_1940(I12887,g4216);
  IV  NOT_1941(g34984,I33252);
  IV  NOT_1942(g32615,g31376);
  IV  NOT_1943(I15834,g11164);
  IV  NOT_1944(g13209,g10632);
  IV  NOT_1945(g8848,g358);
  IV  NOT_1946(g20213,g17062);
  IV  NOT_1947(I15208,g637);
  IV  NOT_1948(g33917,I31779);
  IV  NOT_1949(g21184,g15509);
  IV  NOT_1950(g34419,g34151);
  IV  NOT_1951(g9615,I13236);
  IV  NOT_1952(g21674,g16540);
  IV  NOT_1953(g10812,I14050);
  IV  NOT_1954(g32720,g31710);
  IV  NOT_1955(g30155,I28390);
  IV  NOT_1956(g8398,I12563);
  IV  NOT_1957(g28325,g27463);
  IV  NOT_1958(g12779,g9444);
  IV  NOT_1959(g22898,g20283);
  IV  NOT_1960(g9174,g1205);
  IV  NOT_1961(g34418,g34150);
  IV  NOT_1962(g17794,g13350);
  IV  NOT_1963(g26836,g24866);
  IV  NOT_1964(g17845,I18835);
  IV  NOT_1965(g9374,g5188);
  IV  NOT_1966(g20574,g17847);
  IV  NOT_1967(g20452,g17200);
  IV  NOT_1968(I15542,g1570);
  IV  NOT_1969(g32430,g30984);
  IV  NOT_1970(g10033,g655);
  IV  NOT_1971(g10371,g6918);
  IV  NOT_1972(g32746,g30735);
  IV  NOT_1973(g32493,g30735);
  IV  NOT_1974(g22719,I22024);
  IV  NOT_1975(g24452,g22722);
  IV  NOT_1976(I26100,g26365);
  IV  NOT_1977(g7936,g1061);
  IV  NOT_1978(g9985,g4332);
  IV  NOT_1979(g24047,g19919);
  IV  NOT_1980(g12778,g9856);
  IV  NOT_1981(I18245,g14676);
  IV  NOT_1982(I12764,g4194);
  IV  NOT_1983(g23732,g18833);
  IV  NOT_1984(g8241,g1792);
  IV  NOT_1985(I20793,g17694);
  IV  NOT_1986(g20912,g15171);
  IV  NOT_1987(g19602,g16349);
  IV  NOT_1988(g32465,g30825);
  IV  NOT_1989(g7117,I11816);
  IV  NOT_1990(I18323,g13680);
  IV  NOT_1991(g19657,g16349);
  IV  NOT_1992(g22718,g20887);
  IV  NOT_1993(g16740,g13980);
  IV  NOT_1994(I12132,g577);
  IV  NOT_1995(g19068,g16031);
  IV  NOT_1996(g15169,I17094);
  IV  NOT_1997(g28121,g27093);
  IV  NOT_1998(g9284,g2161);
  IV  NOT_1999(g19375,I19863);
  IV  NOT_2000(g10795,g7202);
  IV  NOT_2001(I25692,g25689);
  IV  NOT_2002(g9239,g5511);
  IV  NOT_2003(g33923,I31791);
  IV  NOT_2004(g9180,g3719);
  IV  NOT_2005(g16186,g13555);
  IV  NOT_2006(g16676,I17876);
  IV  NOT_2007(g16685,g14038);
  IV  NOT_2008(I20690,g15733);
  IV  NOT_2009(I29936,g30606);
  IV  NOT_2010(I17658,g13394);
  IV  NOT_2011(g9380,g5471);
  IV  NOT_2012(g12945,g12467);
  IV  NOT_2013(g31624,I29218);
  IV  NOT_2014(g32806,g31710);
  IV  NOT_2015(g20072,g17384);
  IV  NOT_2016(g32684,g30673);
  IV  NOT_2017(g33688,I31523);
  IV  NOT_2018(g29707,g28504);
  IV  NOT_2019(g9832,g2399);
  IV  NOT_2020(I15073,g10109);
  IV  NOT_2021(g19878,g17271);
  IV  NOT_2022(g24051,g21127);
  IV  NOT_2023(g24072,g20982);
  IV  NOT_2024(g34589,I32675);
  IV  NOT_2025(g17718,g14776);
  IV  NOT_2026(g17521,g14727);
  IV  NOT_2027(g16654,g14136);
  IV  NOT_2028(g20592,g15277);
  IV  NOT_2029(g27998,I26512);
  IV  NOT_2030(I16575,g3298);
  IV  NOT_2031(g15479,g14895);
  IV  NOT_2032(g9853,g5297);
  IV  NOT_2033(I15593,g11989);
  IV  NOT_2034(g8644,g3352);
  IV  NOT_2035(g6989,g4575);
  IV  NOT_2036(g9020,g4287);
  IV  NOT_2037(g24756,g22763);
  IV  NOT_2038(I32452,g34241);
  IV  NOT_2039(I12709,g4284);
  IV  NOT_2040(g21400,g17847);
  IV  NOT_2041(g20780,g15509);
  IV  NOT_2042(g7922,g1312);
  IV  NOT_2043(g8119,g3727);
  IV  NOT_2044(g13530,g12641);
  IV  NOT_2045(g23400,g20676);
  IV  NOT_2046(g12998,g11829);
  IV  NOT_2047(g34836,I33050);
  IV  NOT_2048(g13593,g10556);
  IV  NOT_2049(g28173,I26693);
  IV  NOT_2050(g18929,g16100);
  IV  NOT_2051(g32517,g31194);
  IV  NOT_2052(g23013,g20330);
  IV  NOT_2053(I28572,g28274);
  IV  NOT_2054(g12233,g10338);
  IV  NOT_2055(I31586,g33149);
  IV  NOT_2056(g23214,g20785);
  IV  NOT_2057(g11122,g8751);
  IV  NOT_2058(I14902,g9821);
  IV  NOT_2059(I14301,g8571);
  IV  NOT_2060(g12182,I15030);
  IV  NOT_2061(g29978,g28927);
  IV  NOT_2062(g12672,g10003);
  IV  NOT_2063(g7581,g1379);
  IV  NOT_2064(g21329,g16577);
  IV  NOT_2065(g22926,g20391);
  IV  NOT_2066(g25155,g22472);
  IV  NOT_2067(g9559,g6077);
  IV  NOT_2068(g13565,g11006);
  IV  NOT_2069(g6971,I11737);
  IV  NOT_2070(g8818,I12808);
  IV  NOT_2071(I25005,g24417);
  IV  NOT_2072(g14421,I16575);
  IV  NOT_2073(I19704,g17653);
  IV  NOT_2074(g25266,g22228);
  IV  NOT_2075(g25170,g22498);
  IV  NOT_2076(g9931,g5763);
  IV  NOT_2077(g23539,g21070);
  IV  NOT_2078(g17573,g12911);
  IV  NOT_2079(g7597,g952);
  IV  NOT_2080(g11034,g7611);
  IV  NOT_2081(g23005,g20283);
  IV  NOT_2082(g13034,g11920);
  IV  NOT_2083(g17247,I18259);
  IV  NOT_2084(I32051,g33631);
  IV  NOT_2085(g30022,g29001);
  IV  NOT_2086(g34118,I32051);
  IV  NOT_2087(I16606,g3649);
  IV  NOT_2088(g15580,g13242);
  IV  NOT_2089(g12932,I15550);
  IV  NOT_2090(g23538,g20924);
  IV  NOT_2091(g34864,g34840);
  IV  NOT_2092(I16492,g12430);
  IV  NOT_2093(g17389,g14915);
  IV  NOT_2094(g17926,I18852);
  IV  NOT_2095(g16964,I18120);
  IV  NOT_2096(g24152,I23300);
  IV  NOT_2097(g19458,I19927);
  IV  NOT_2098(g30313,g28843);
  IV  NOT_2099(g34749,I32921);
  IV  NOT_2100(g17612,g15014);
  IV  NOT_2101(g24396,g22885);
  IV  NOT_2102(g8211,g2319);
  IV  NOT_2103(g29067,I27401);
  IV  NOT_2104(g9905,g802);
  IV  NOT_2105(g10541,g9407);
  IV  NOT_2106(g16423,g14066);
  IV  NOT_2107(g27961,g26816);
  IV  NOT_2108(g8186,g990);
  IV  NOT_2109(g34313,g34086);
  IV  NOT_2110(I13552,g121);
  IV  NOT_2111(g10473,I13857);
  IV  NOT_2112(g17324,I18301);
  IV  NOT_2113(g32523,g30825);
  IV  NOT_2114(I24128,g23009);
  IV  NOT_2115(g31854,g29385);
  IV  NOT_2116(g14541,g11405);
  IV  NOT_2117(g16216,I17557);
  IV  NOT_2118(I29909,g31791);
  IV  NOT_2119(I33041,g34772);
  IV  NOT_2120(g12897,g10400);
  IV  NOT_2121(g13409,I15918);
  IV  NOT_2122(g16587,I17763);
  IV  NOT_2123(g17777,g14908);
  IV  NOT_2124(g25167,I24331);
  IV  NOT_2125(g25194,g22763);
  IV  NOT_2126(I13779,g6868);
  IV  NOT_2127(I26584,g26943);
  IV  NOT_2128(g9630,g6527);
  IV  NOT_2129(g29150,g27886);
  IV  NOT_2130(g34276,g34058);
  IV  NOT_2131(g34285,I32284);
  IV  NOT_2132(g7995,g153);
  IV  NOT_2133(g30305,g28939);
  IV  NOT_2134(g11136,I14192);
  IV  NOT_2135(g30053,g29121);
  IV  NOT_2136(g8026,g3857);
  IV  NOT_2137(g25524,g22228);
  IV  NOT_2138(I27970,g28803);
  IV  NOT_2139(g18827,g16000);
  IV  NOT_2140(g34053,g33683);
  IV  NOT_2141(g7479,g1008);
  IV  NOT_2142(g9300,g5180);
  IV  NOT_2143(g10359,g6830);
  IV  NOT_2144(I32820,g34474);
  IV  NOT_2145(g8426,g3045);
  IV  NOT_2146(g32475,g30614);
  IV  NOT_2147(g14359,I16515);
  IV  NOT_2148(g8170,g3770);
  IV  NOT_2149(g7840,g4878);
  IV  NOT_2150(g22997,g20391);
  IV  NOT_2151(g32727,g31710);
  IV  NOT_2152(g10358,g6827);
  IV  NOT_2153(g33660,I31494);
  IV  NOT_2154(g32863,g31021);
  IV  NOT_2155(g29196,g27059);
  IV  NOT_2156(I32846,g34502);
  IV  NOT_2157(g14535,g12318);
  IV  NOT_2158(g24405,g22722);
  IV  NOT_2159(g8125,g3869);
  IV  NOT_2160(g30036,g29085);
  IV  NOT_2161(g14358,I16512);
  IV  NOT_2162(g25119,g22384);
  IV  NOT_2163(I22819,g19862);
  IV  NOT_2164(g8821,I12811);
  IV  NOT_2165(g16000,I17425);
  IV  NOT_2166(g15740,g13342);
  IV  NOT_2167(I25683,g25642);
  IV  NOT_2168(I29242,g29313);
  IV  NOT_2169(g32437,I29965);
  IV  NOT_2170(g14828,I16875);
  IV  NOT_2171(g23235,g20785);
  IV  NOT_2172(g33456,I30986);
  IV  NOT_2173(g10121,g2327);
  IV  NOT_2174(g11164,g8085);
  IV  NOT_2175(g25118,g22417);
  IV  NOT_2176(g26693,g25300);
  IV  NOT_2177(g8280,g3443);
  IV  NOT_2178(g23683,I22816);
  IV  NOT_2179(g15373,I17118);
  IV  NOT_2180(g9973,g2112);
  IV  NOT_2181(g33916,I31776);
  IV  NOT_2182(I22111,g19919);
  IV  NOT_2183(g7356,g1802);
  IV  NOT_2184(I17819,g3618);
  IV  NOT_2185(g16747,g14113);
  IV  NOT_2186(g20583,g17873);
  IV  NOT_2187(g32703,g30825);
  IV  NOT_2188(I12994,g6748);
  IV  NOT_2189(I15474,g10364);
  IV  NOT_2190(g24020,g20014);
  IV  NOT_2191(g19532,g16821);
  IV  NOT_2192(g22360,I21849);
  IV  NOT_2193(g9040,g499);
  IV  NOT_2194(g28648,g27693);
  IV  NOT_2195(g18881,I19671);
  IV  NOT_2196(I13672,g106);
  IV  NOT_2197(g13474,g11048);
  IV  NOT_2198(I25882,g25776);
  IV  NOT_2199(g20046,g16540);
  IV  NOT_2200(g9969,g1682);
  IV  NOT_2201(g19783,g16931);
  IV  NOT_2202(I17111,g13809);
  IV  NOT_2203(g16123,g13530);
  IV  NOT_2204(g24046,g21256);
  IV  NOT_2205(g17871,I18845);
  IV  NOT_2206(g16814,g14058);
  IV  NOT_2207(g21414,g17929);
  IV  NOT_2208(g32600,g31542);
  IV  NOT_2209(g7704,I12167);
  IV  NOT_2210(I16663,g10981);
  IV  NOT_2211(g23515,g20785);
  IV  NOT_2212(g28604,g27759);
  IV  NOT_2213(g23882,g19277);
  IV  NOT_2214(g23414,I22525);
  IV  NOT_2215(g32781,g31376);
  IV  NOT_2216(I23099,g20682);
  IV  NOT_2217(g31596,I29204);
  IV  NOT_2218(g8106,g3133);
  IV  NOT_2219(g14173,g12076);
  IV  NOT_2220(I23324,g21697);
  IV  NOT_2221(g20113,g16826);
  IV  NOT_2222(g21407,g15171);
  IV  NOT_2223(g31243,g29933);
  IV  NOT_2224(I17590,g14591);
  IV  NOT_2225(g19353,I19831);
  IV  NOT_2226(g24113,g19984);
  IV  NOT_2227(I32929,g34649);
  IV  NOT_2228(g32952,g30937);
  IV  NOT_2229(g19144,g16031);
  IV  NOT_2230(g12811,g10319);
  IV  NOT_2231(g27971,g26673);
  IV  NOT_2232(g8187,g1657);
  IV  NOT_2233(g32821,g31021);
  IV  NOT_2234(g8387,g3080);
  IV  NOT_2235(g25036,g23733);
  IV  NOT_2236(I31523,g33187);
  IV  NOT_2237(g7163,g4593);
  IV  NOT_2238(g29597,g28444);
  IV  NOT_2239(g25101,g22384);
  IV  NOT_2240(g20105,g17433);
  IV  NOT_2241(g24357,g22325);
  IV  NOT_2242(g25560,g22550);
  IV  NOT_2243(g10029,I13548);
  IV  NOT_2244(g8756,g4049);
  IV  NOT_2245(g22220,I21802);
  IV  NOT_2246(g13303,I15869);
  IV  NOT_2247(g24105,g19935);
  IV  NOT_2248(I17094,g14331);
  IV  NOT_2249(I18031,g13680);
  IV  NOT_2250(g29689,I27954);
  IV  NOT_2251(g14029,g11283);
  IV  NOT_2252(g29923,g28874);
  IV  NOT_2253(g25642,I24787);
  IV  NOT_2254(g32790,g30825);
  IV  NOT_2255(g9648,g2177);
  IV  NOT_2256(g32137,g31134);
  IV  NOT_2257(g10028,g8);
  IV  NOT_2258(g9875,g5747);
  IV  NOT_2259(g32516,g31070);
  IV  NOT_2260(g31655,I29233);
  IV  NOT_2261(I29579,g30565);
  IV  NOT_2262(g28262,I26785);
  IV  NOT_2263(I24445,g22923);
  IV  NOT_2264(g20640,g15426);
  IV  NOT_2265(I17801,g14936);
  IV  NOT_2266(g20769,g17955);
  IV  NOT_2267(g17472,g14656);
  IV  NOT_2268(I26406,g26187);
  IV  NOT_2269(g12368,I15208);
  IV  NOT_2270(I16040,g10430);
  IV  NOT_2271(I20499,g16224);
  IV  NOT_2272(I12086,g622);
  IV  NOT_2273(g33670,I31504);
  IV  NOT_2274(I31727,g33076);
  IV  NOT_2275(g32873,g30614);
  IV  NOT_2276(g8046,g528);
  IV  NOT_2277(g25064,I24228);
  IV  NOT_2278(g16510,g14008);
  IV  NOT_2279(g19364,g15825);
  IV  NOT_2280(g20768,g17955);
  IV  NOT_2281(g28633,g27687);
  IV  NOT_2282(g8514,g4258);
  IV  NOT_2283(I19238,g15079);
  IV  NOT_2284(g34570,g34392);
  IV  NOT_2285(g34712,I32868);
  IV  NOT_2286(g21725,I21294);
  IV  NOT_2287(g11796,g7985);
  IV  NOT_2288(g16579,g13267);
  IV  NOT_2289(g33335,I30861);
  IV  NOT_2290(g8403,I12568);
  IV  NOT_2291(g23759,I22886);
  IV  NOT_2292(g13174,g10741);
  IV  NOT_2293(I21766,g19620);
  IV  NOT_2294(I17695,g14330);
  IV  NOT_2295(g26941,I25689);
  IV  NOT_2296(g34914,I33134);
  IV  NOT_2297(g31839,g29385);
  IV  NOT_2298(g33839,I31686);
  IV  NOT_2299(I32827,g34477);
  IV  NOT_2300(g8345,g3794);
  IV  NOT_2301(g8841,I12823);
  IV  NOT_2302(I14671,g7717);
  IV  NOT_2303(g7157,g5706);
  IV  NOT_2304(I12159,g608);
  IV  NOT_2305(g22147,g18997);
  IV  NOT_2306(g26519,I25380);
  IV  NOT_2307(g16578,I17750);
  IV  NOT_2308(g15569,I17148);
  IV  NOT_2309(g8763,I12749);
  IV  NOT_2310(I16564,g10429);
  IV  NOT_2311(g23435,g18833);
  IV  NOT_2312(g31667,g30142);
  IV  NOT_2313(g31838,g29385);
  IV  NOT_2314(g23082,g21024);
  IV  NOT_2315(g32834,g31672);
  IV  NOT_2316(g9839,g2724);
  IV  NOT_2317(g30074,g29046);
  IV  NOT_2318(g26518,g25233);
  IV  NOT_2319(g17591,I18526);
  IV  NOT_2320(g12896,g10402);
  IV  NOT_2321(g17776,g14905);
  IV  NOT_2322(g27011,g25917);
  IV  NOT_2323(I27561,g28163);
  IV  NOT_2324(g15568,g14984);
  IV  NOT_2325(g15747,g13307);
  IV  NOT_2326(g25009,g22472);
  IV  NOT_2327(I13723,g3167);
  IV  NOT_2328(I26004,g26818);
  IV  NOT_2329(I18868,g14315);
  IV  NOT_2330(I23360,g23360);
  IV  NOT_2331(g18945,g16100);
  IV  NOT_2332(g30567,g29930);
  IV  NOT_2333(I30962,g32021);
  IV  NOT_2334(g17147,g14321);
  IV  NOT_2335(g22858,g20751);
  IV  NOT_2336(g34594,I32690);
  IV  NOT_2337(I13149,g6745);
  IV  NOT_2338(g17754,g14262);
  IV  NOT_2339(I16847,g6329);
  IV  NOT_2340(g26935,I25677);
  IV  NOT_2341(g25008,g22432);
  IV  NOT_2342(g32542,g31554);
  IV  NOT_2343(g8107,g3179);
  IV  NOT_2344(I32803,g34584);
  IV  NOT_2345(I25399,g24489);
  IV  NOT_2346(g31487,I29149);
  IV  NOT_2347(g32021,I29579);
  IV  NOT_2348(g32453,I29981);
  IV  NOT_2349(I29720,g30931);
  IV  NOT_2350(g11192,g8038);
  IV  NOT_2351(g22151,I21734);
  IV  NOT_2352(I11620,g1);
  IV  NOT_2353(I21162,g17292);
  IV  NOT_2354(I12144,g554);
  IV  NOT_2355(I12823,g4311);
  IV  NOT_2356(I18709,g6668);
  IV  NOT_2357(g20662,g15171);
  IV  NOT_2358(g21399,g15224);
  IV  NOT_2359(g23849,g19277);
  IV  NOT_2360(g22996,g20330);
  IV  NOT_2361(g23940,g19074);
  IV  NOT_2362(g25892,g24528);
  IV  NOT_2363(I20753,g16677);
  IV  NOT_2364(I15663,g5308);
  IV  NOT_2365(g23399,g21514);
  IV  NOT_2366(g32726,g31672);
  IV  NOT_2367(g32913,g30825);
  IV  NOT_2368(g24027,g20014);
  IV  NOT_2369(I18259,g12946);
  IV  NOT_2370(g9618,g5794);
  IV  NOT_2371(g11663,g6905);
  IV  NOT_2372(g16615,I17801);
  IV  NOT_2373(g22844,g21163);
  IV  NOT_2374(g13522,g10981);
  IV  NOT_2375(g34941,g34926);
  IV  NOT_2376(g13663,g10971);
  IV  NOT_2377(g21398,g18008);
  IV  NOT_2378(g23848,g19210);
  IV  NOT_2379(g25555,g22550);
  IV  NOT_2380(g32614,g31542);
  IV  NOT_2381(g7626,I12112);
  IV  NOT_2382(I12336,g52);
  IV  NOT_2383(g23398,g21468);
  IV  NOT_2384(I32881,g34688);
  IV  NOT_2385(g8858,g671);
  IV  NOT_2386(g33443,I30971);
  IV  NOT_2387(g16720,g14234);
  IV  NOT_2388(g9282,g723);
  IV  NOT_2389(g34675,I32809);
  IV  NOT_2390(I20650,g17010);
  IV  NOT_2391(g23652,I22785);
  IV  NOT_2392(g32607,g31542);
  IV  NOT_2393(g8016,g3391);
  IV  NOT_2394(g10981,I14119);
  IV  NOT_2395(g8757,I12746);
  IV  NOT_2396(g32905,g30825);
  IV  NOT_2397(g14563,I16676);
  IV  NOT_2398(g8416,I12580);
  IV  NOT_2399(g27112,g26793);
  IV  NOT_2400(g20710,g15509);
  IV  NOT_2401(g16746,g14258);
  IV  NOT_2402(I20529,g16309);
  IV  NOT_2403(I21911,g21278);
  IV  NOT_2404(g17844,I18832);
  IV  NOT_2405(g20552,g17847);
  IV  NOT_2406(g32530,g30825);
  IV  NOT_2407(g9693,g1886);
  IV  NOT_2408(g13483,g11270);
  IV  NOT_2409(I33264,g34978);
  IV  NOT_2410(I15862,g11215);
  IV  NOT_2411(g17367,I18320);
  IV  NOT_2412(g32593,g31542);
  IV  NOT_2413(g18932,g16136);
  IV  NOT_2414(g6985,g4669);
  IV  NOT_2415(I33137,g34884);
  IV  NOT_2416(g20204,g16578);
  IV  NOT_2417(g19687,g17096);
  IV  NOT_2418(I21246,g16540);
  IV  NOT_2419(g24003,g21514);
  IV  NOT_2420(g23263,I22366);
  IV  NOT_2421(I12631,g1242);
  IV  NOT_2422(g8522,g298);
  IV  NOT_2423(g20779,g15509);
  IV  NOT_2424(g22319,I21831);
  IV  NOT_2425(g12378,g9417);
  IV  NOT_2426(g34935,I33189);
  IV  NOT_2427(g23332,g20785);
  IV  NOT_2428(g32565,g30735);
  IV  NOT_2429(g32464,g30735);
  IV  NOT_2430(g25239,g23972);
  IV  NOT_2431(g19954,g16540);
  IV  NOT_2432(g11949,I14773);
  IV  NOT_2433(I24393,g23453);
  IV  NOT_2434(g19374,g16047);
  IV  NOT_2435(g20778,g15224);
  IV  NOT_2436(g34883,g34852);
  IV  NOT_2437(g10794,g8470);
  IV  NOT_2438(g9555,I13206);
  IV  NOT_2439(g18897,g15509);
  IV  NOT_2440(I15536,g1227);
  IV  NOT_2441(g10395,g6995);
  IV  NOT_2442(g22227,g19801);
  IV  NOT_2443(g24778,g23286);
  IV  NOT_2444(g9804,g5456);
  IV  NOT_2445(g10262,g586);
  IV  NOT_2446(g24081,g21209);
  IV  NOT_2447(g21406,g17955);
  IV  NOT_2448(g16684,g14223);
  IV  NOT_2449(g11948,g10224);
  IV  NOT_2450(I21776,g21308);
  IV  NOT_2451(I15702,g12217);
  IV  NOT_2452(g14262,g10838);
  IV  NOT_2453(g12944,g12659);
  IV  NOT_2454(I18810,g13716);
  IV  NOT_2455(g23406,g20330);
  IV  NOT_2456(g9792,g5401);
  IV  NOT_2457(g32641,g30614);
  IV  NOT_2458(g6832,I11665);
  IV  NOT_2459(g32797,g30825);
  IV  NOT_2460(g23962,g19147);
  IV  NOT_2461(g31815,g29385);
  IV  NOT_2462(g23361,I22464);
  IV  NOT_2463(g28032,g26365);
  IV  NOT_2464(I32482,g34304);
  IV  NOT_2465(g11702,g6928);
  IV  NOT_2466(g7778,g1339);
  IV  NOT_2467(g15579,I17159);
  IV  NOT_2468(g31601,I29207);
  IV  NOT_2469(g8654,g1087);
  IV  NOT_2470(I16452,g11182);
  IV  NOT_2471(I18879,g13267);
  IV  NOT_2472(g9621,g6423);
  IV  NOT_2473(g10191,g6386);
  IV  NOT_2474(g23500,g20924);
  IV  NOT_2475(g24356,g22594);
  IV  NOT_2476(g13621,g10573);
  IV  NOT_2477(g21049,g17433);
  IV  NOT_2478(I11896,g4446);
  IV  NOT_2479(g25185,g22228);
  IV  NOT_2480(g17059,I18151);
  IV  NOT_2481(g20380,g17955);
  IV  NOT_2482(g26083,g24809);
  IV  NOT_2483(g14191,g12381);
  IV  NOT_2484(g30729,I28883);
  IV  NOT_2485(I15564,g11949);
  IV  NOT_2486(g25092,g23666);
  IV  NOT_2487(g24999,g23626);
  IV  NOT_2488(g26284,g24875);
  IV  NOT_2489(I18337,g1422);
  IV  NOT_2490(g34501,g34400);
  IV  NOT_2491(g27730,g26424);
  IV  NOT_2492(g10521,I13889);
  IV  NOT_2493(g12857,I15474);
  IV  NOT_2494(I19348,g15084);
  IV  NOT_2495(g21048,g17533);
  IV  NOT_2496(g25154,g22457);
  IV  NOT_2497(g20090,g17433);
  IV  NOT_2498(g17058,I18148);
  IV  NOT_2499(g32635,g31542);
  IV  NOT_2500(g8880,I12861);
  IV  NOT_2501(g31937,g30991);
  IV  NOT_2502(g8595,I12666);
  IV  NOT_2503(g24090,g19935);
  IV  NOT_2504(g19489,g16449);
  IV  NOT_2505(g20233,g17873);
  IV  NOT_2506(g33937,I31823);
  IV  NOT_2507(g12793,g10287);
  IV  NOT_2508(I11716,g4054);
  IV  NOT_2509(g20182,g16897);
  IV  NOT_2510(g20651,g15483);
  IV  NOT_2511(g20672,g15277);
  IV  NOT_2512(I17876,g13070);
  IV  NOT_2513(g23004,g20283);
  IV  NOT_2514(I27495,g27961);
  IV  NOT_2515(g7475,g896);
  IV  NOT_2516(g21221,g15680);
  IV  NOT_2517(g24182,I23390);
  IV  NOT_2518(g19559,g16129);
  IV  NOT_2519(g23221,g20785);
  IV  NOT_2520(I14644,g7717);
  IV  NOT_2521(g11183,g8135);
  IV  NOT_2522(g29942,g28867);
  IV  NOT_2523(g22957,I22143);
  IV  NOT_2524(g31791,I29363);
  IV  NOT_2525(g7627,g4311);
  IV  NOT_2526(g19558,g15938);
  IV  NOT_2527(g6905,I11708);
  IV  NOT_2528(g16523,g14041);
  IV  NOT_2529(g8612,g2775);
  IV  NOT_2530(g23613,I22748);
  IV  NOT_2531(g9518,g6219);
  IV  NOT_2532(g15615,I17181);
  IV  NOT_2533(I17763,g13191);
  IV  NOT_2534(I31607,g33164);
  IV  NOT_2535(g13062,g10981);
  IV  NOT_2536(g7526,I12013);
  IV  NOT_2537(g7998,g392);
  IV  NOT_2538(g11509,g7632);
  IV  NOT_2539(g22146,g18997);
  IV  NOT_2540(g26653,g25337);
  IV  NOT_2541(g20513,g18065);
  IV  NOT_2542(g17301,g14454);
  IV  NOT_2543(g20449,g15277);
  IV  NOT_2544(g28162,I26679);
  IV  NOT_2545(g10389,g6986);
  IV  NOT_2546(g32891,g30825);
  IV  NOT_2547(I15872,g11236);
  IV  NOT_2548(g13933,g11419);
  IV  NOT_2549(g23947,g19210);
  IV  NOT_2550(g31479,I29139);
  IV  NOT_2551(g31666,I29248);
  IV  NOT_2552(I27954,g28803);
  IV  NOT_2553(g18097,I18897);
  IV  NOT_2554(g21273,I21006);
  IV  NOT_2555(g17120,g14262);
  IV  NOT_2556(g19544,g16349);
  IV  NOT_2557(g23273,g21070);
  IV  NOT_2558(g19865,g15885);
  IV  NOT_2559(g17739,I18728);
  IV  NOT_2560(g10612,g10233);
  IV  NOT_2561(g11872,I14684);
  IV  NOT_2562(g23605,g20739);
  IV  NOT_2563(g9776,g5073);
  IV  NOT_2564(g10099,g6682);
  IV  NOT_2565(g15746,g13121);
  IV  NOT_2566(g16475,g14107);
  IV  NOT_2567(g20448,g15509);
  IV  NOT_2568(g34304,I32309);
  IV  NOT_2569(I12954,g4358);
  IV  NOT_2570(g10388,g6983);
  IV  NOT_2571(I32651,g34375);
  IV  NOT_2572(g32575,g31170);
  IV  NOT_2573(g32474,g31194);
  IV  NOT_2574(g19713,g16816);
  IV  NOT_2575(g7439,g6351);
  IV  NOT_2576(g29930,I28162);
  IV  NOT_2577(g22698,I22009);
  IV  NOT_2578(g29993,g29018);
  IV  NOT_2579(g16727,g14454);
  IV  NOT_2580(g17738,g14813);
  IV  NOT_2581(g17645,g15018);
  IV  NOT_2582(g20505,g15426);
  IV  NOT_2583(g21463,g15588);
  IV  NOT_2584(g23812,g18997);
  IV  NOT_2585(g32711,g31070);
  IV  NOT_2586(g8130,g4515);
  IV  NOT_2587(g14701,g12351);
  IV  NOT_2588(I17456,g13680);
  IV  NOT_2589(I23318,g21689);
  IV  NOT_2590(g8542,I12644);
  IV  NOT_2591(g24505,g22689);
  IV  NOT_2592(g8330,g2587);
  IV  NOT_2593(g24404,g22908);
  IV  NOT_2594(g10272,I13705);
  IV  NOT_2595(g9965,g127);
  IV  NOT_2596(g29965,g28903);
  IV  NOT_2597(I33034,g34769);
  IV  NOT_2598(g14251,g12308);
  IV  NOT_2599(I17916,g13087);
  IV  NOT_2600(g20026,g17271);
  IV  NOT_2601(g32537,g30825);
  IV  NOT_2602(I18078,g13350);
  IV  NOT_2603(g20212,g17194);
  IV  NOT_2604(g23234,g20375);
  IV  NOT_2605(g24026,g19919);
  IV  NOT_2606(g9264,g5396);
  IV  NOT_2607(g15806,I17302);
  IV  NOT_2608(I21058,g17747);
  IV  NOT_2609(g25438,g22763);
  IV  NOT_2610(g6973,I11743);
  IV  NOT_2611(I17314,g14078);
  IV  NOT_2612(I32449,g34127);
  IV  NOT_2613(g19679,g16782);
  IV  NOT_2614(I18086,g13856);
  IV  NOT_2615(g27245,g26209);
  IV  NOT_2616(g34653,I32763);
  IV  NOT_2617(g9360,g3372);
  IV  NOT_2618(g9933,g5759);
  IV  NOT_2619(g32606,g30673);
  IV  NOT_2620(g10032,g562);
  IV  NOT_2621(I29236,g29498);
  IV  NOT_2622(g32492,g31376);
  IV  NOT_2623(g19678,g16752);
  IV  NOT_2624(I15205,g10139);
  IV  NOT_2625(g14032,g11048);
  IV  NOT_2626(g10140,g19);
  IV  NOT_2627(g29210,I27546);
  IV  NOT_2628(g9050,g1087);
  IV  NOT_2629(g17427,I18364);
  IV  NOT_2630(I13802,g6971);
  IV  NOT_2631(g13574,I16024);
  IV  NOT_2632(I25514,g25073);
  IV  NOT_2633(I13857,g9780);
  IV  NOT_2634(g17366,g14454);
  IV  NOT_2635(g7952,g3774);
  IV  NOT_2636(g25083,g23782);
  IV  NOT_2637(g25348,g22763);
  IV  NOT_2638(g9450,g5817);
  IV  NOT_2639(I14450,g4191);
  IV  NOT_2640(g16600,I17780);
  IV  NOT_2641(g19686,g17062);
  IV  NOT_2642(g25284,I24474);
  IV  NOT_2643(g21514,I21189);
  IV  NOT_2644(I11793,g6049);
  IV  NOT_2645(g11912,g8989);
  IV  NOT_2646(g26576,I25399);
  IV  NOT_2647(I26682,g27774);
  IV  NOT_2648(g28147,I26654);
  IV  NOT_2649(I27558,g28155);
  IV  NOT_2650(g32750,g30937);
  IV  NOT_2651(I12016,g772);
  IV  NOT_2652(I18125,g13191);
  IV  NOT_2653(g10061,I13581);
  IV  NOT_2654(g13311,I15878);
  IV  NOT_2655(g28754,I27238);
  IV  NOT_2656(g32381,I29909);
  IV  NOT_2657(g7616,I12086);
  IV  NOT_2658(I19484,g15122);
  IV  NOT_2659(g23507,g21562);
  IV  NOT_2660(g34852,g34845);
  IV  NOT_2661(g20433,g17929);
  IV  NOT_2662(g25566,g22550);
  IV  NOT_2663(g18896,g16031);
  IV  NOT_2664(g24149,g19338);
  IV  NOT_2665(g20387,g15426);
  IV  NOT_2666(g28370,g27528);
  IV  NOT_2667(I28866,g29730);
  IV  NOT_2668(I22180,g21366);
  IV  NOT_2669(g16821,I18031);
  IV  NOT_2670(g21421,g15171);
  IV  NOT_2671(g27737,g26718);
  IV  NOT_2672(I12893,g4226);
  IV  NOT_2673(g7004,I11777);
  IV  NOT_2674(g9379,g5424);
  IV  NOT_2675(g23421,g21562);
  IV  NOT_2676(g13051,g11964);
  IV  NOT_2677(g20097,g17691);
  IV  NOT_2678(g32796,g31376);
  IV  NOT_2679(g7527,I12016);
  IV  NOT_2680(I33164,g34894);
  IV  NOT_2681(g24097,g19935);
  IV  NOT_2682(g26608,g25334);
  IV  NOT_2683(g11592,I14537);
  IV  NOT_2684(g20104,g17433);
  IV  NOT_2685(g7647,I12132);
  IV  NOT_2686(g34664,I32782);
  IV  NOT_2687(I27713,g28224);
  IV  NOT_2688(I13548,g94);
  IV  NOT_2689(g10360,g6836);
  IV  NOT_2690(g23012,g20330);
  IV  NOT_2691(g24104,g19890);
  IV  NOT_2692(g17226,I18252);
  IV  NOT_2693(g25139,g22472);
  IV  NOT_2694(g17715,I18700);
  IV  NOT_2695(g6875,I11697);
  IV  NOT_2696(g9777,g5112);
  IV  NOT_2697(g17481,g15005);
  IV  NOT_2698(I25541,g25180);
  IV  NOT_2699(g32840,g30825);
  IV  NOT_2700(I28597,g29374);
  IV  NOT_2701(g28367,I26880);
  IV  NOT_2702(I31474,g33212);
  IV  NOT_2703(g24971,g23590);
  IV  NOT_2704(g27880,I26427);
  IV  NOT_2705(g25138,g22472);
  IV  NOT_2706(g34576,I32654);
  IV  NOT_2707(g16873,I18063);
  IV  NOT_2708(g23541,g21514);
  IV  NOT_2709(g31800,g29385);
  IV  NOT_2710(g12995,g11820);
  IV  NOT_2711(g7503,g1351);
  IV  NOT_2712(g7970,g4688);
  IV  NOT_2713(g13350,I15906);
  IV  NOT_2714(g23473,g20785);
  IV  NOT_2715(g33800,I31642);
  IV  NOT_2716(g8056,g1246);
  IV  NOT_2717(I13317,g6144);
  IV  NOT_2718(g11820,I14644);
  IV  NOT_2719(g33936,I31820);
  IV  NOT_2720(g8456,g56);
  IV  NOT_2721(g12880,g10387);
  IV  NOT_2722(I22131,g19984);
  IV  NOT_2723(I24078,g22360);
  IV  NOT_2724(g23789,g21308);
  IV  NOT_2725(I17839,g13412);
  IV  NOT_2726(g32192,g31262);
  IV  NOT_2727(I33109,g34851);
  IV  NOT_2728(I15846,g11183);
  IV  NOT_2729(I16357,g884);
  IV  NOT_2730(I25359,g24715);
  IV  NOT_2731(I19799,g17817);
  IV  NOT_2732(g30312,g28970);
  IV  NOT_2733(I12189,g5869);
  IV  NOT_2734(I19813,g17952);
  IV  NOT_2735(g24368,g22228);
  IV  NOT_2736(g21724,I21291);
  IV  NOT_2737(g23788,g18997);
  IV  NOT_2738(g8155,g3380);
  IV  NOT_2739(g34312,g34098);
  IV  NOT_2740(g26973,g26105);
  IV  NOT_2741(g34200,g33895);
  IV  NOT_2742(g7224,g4601);
  IV  NOT_2743(g32522,g30735);
  IV  NOT_2744(g23359,I22458);
  IV  NOT_2745(g32663,g30673);
  IV  NOT_2746(g8355,I12534);
  IV  NOT_2747(g8851,g590);
  IV  NOT_2748(I13057,g112);
  IV  NOT_2749(g14451,I16606);
  IV  NOT_2750(I23366,g23321);
  IV  NOT_2751(I18364,g13009);
  IV  NOT_2752(I22619,g21193);
  IV  NOT_2753(I17131,g14384);
  IV  NOT_2754(I22502,g19376);
  IV  NOT_2755(g22980,I22153);
  IV  NOT_2756(g21434,g17248);
  IV  NOT_2757(I22557,g20695);
  IV  NOT_2758(g21358,g16307);
  IV  NOT_2759(g6839,g1858);
  IV  NOT_2760(g23434,g21611);
  IV  NOT_2761(g24850,I24022);
  IV  NOT_2762(g30052,g29018);
  IV  NOT_2763(I19674,g15932);
  IV  NOT_2764(g8964,g4269);
  IV  NOT_2765(I29913,g30605);
  IV  NOT_2766(g27831,I26406);
  IV  NOT_2767(I11626,g31);
  IV  NOT_2768(g11413,g9100);
  IV  NOT_2769(g34921,I33155);
  IV  NOT_2770(g13413,g11737);
  IV  NOT_2771(g34052,g33635);
  IV  NOT_2772(g23946,g19210);
  IV  NOT_2773(g24133,g19935);
  IV  NOT_2774(g29169,g27886);
  IV  NOT_2775(g18096,I18894);
  IV  NOT_2776(g18944,g15938);
  IV  NOT_2777(g20229,g17015);
  IV  NOT_2778(g32483,g30673);
  IV  NOT_2779(g19617,g16349);
  IV  NOT_2780(g19470,g16000);
  IV  NOT_2781(g22181,g19277);
  IV  NOT_2782(g11691,I14570);
  IV  NOT_2783(g19915,g16349);
  IV  NOT_2784(g12831,g9569);
  IV  NOT_2785(g26732,g25389);
  IV  NOT_2786(I16803,g6369);
  IV  NOT_2787(I12030,g595);
  IV  NOT_2788(I17557,g14510);
  IV  NOT_2789(g9541,g2012);
  IV  NOT_2790(g32553,g31170);
  IV  NOT_2791(g32862,g30825);
  IV  NOT_2792(g7617,I12089);
  IV  NOT_2793(g16726,g14454);
  IV  NOT_2794(I26649,g27675);
  IV  NOT_2795(g34813,I33027);
  IV  NOT_2796(g10776,I14033);
  IV  NOT_2797(g19277,I19813);
  IV  NOT_2798(g32949,g30825);
  IV  NOT_2799(g9332,g64);
  IV  NOT_2800(g14591,I16709);
  IV  NOT_2801(g14785,g12629);
  IV  NOT_2802(I21226,g16540);
  IV  NOT_2803(I22286,g19446);
  IV  NOT_2804(g7516,I12003);
  IV  NOT_2805(g21682,g16540);
  IV  NOT_2806(I18224,g13793);
  IV  NOT_2807(g9680,I13276);
  IV  NOT_2808(g9153,I12991);
  IV  NOT_2809(g10147,g728);
  IV  NOT_2810(g20716,g15277);
  IV  NOT_2811(g27989,g26759);
  IV  NOT_2812(g29217,I27567);
  IV  NOT_2813(g34973,I33235);
  IV  NOT_2814(g25554,g22550);
  IV  NOT_2815(I15929,g10430);
  IV  NOT_2816(I18571,g13074);
  IV  NOT_2817(g21291,g16620);
  IV  NOT_2818(g32536,g31376);
  IV  NOT_2819(g14147,I16357);
  IV  NOT_2820(g30184,g28144);
  IV  NOT_2821(I31796,g33176);
  IV  NOT_2822(g10355,g6816);
  IV  NOT_2823(g32948,g30735);
  IV  NOT_2824(g23291,g21070);
  IV  NOT_2825(g16607,g13960);
  IV  NOT_2826(g19494,g16349);
  IV  NOT_2827(g11929,I14745);
  IV  NOT_2828(I11737,g4467);
  IV  NOT_2829(g34674,I32806);
  IV  NOT_2830(g8279,I12487);
  IV  NOT_2831(g16320,g14454);
  IV  NOT_2832(g20582,g17873);
  IV  NOT_2833(g32702,g30735);
  IV  NOT_2834(g9744,g6486);
  IV  NOT_2835(g10370,g7095);
  IV  NOT_2836(g31000,g29737);
  IV  NOT_2837(g32757,g30937);
  IV  NOT_2838(g32904,g30735);
  IV  NOT_2839(g6988,g4765);
  IV  NOT_2840(I14866,g9748);
  IV  NOT_2841(g16530,g14454);
  IV  NOT_2842(g26400,I25351);
  IV  NOT_2843(g11928,I14742);
  IV  NOT_2844(g25115,I24281);
  IV  NOT_2845(g13583,I16028);
  IV  NOT_2846(g32621,g31542);
  IV  NOT_2847(g8872,g4258);
  IV  NOT_2848(g22520,g19801);
  IV  NOT_2849(I22601,g21127);
  IV  NOT_2850(g10151,g1992);
  IV  NOT_2851(g28120,g27108);
  IV  NOT_2852(I32228,g34122);
  IV  NOT_2853(I11697,g3352);
  IV  NOT_2854(g10172,g6459);
  IV  NOT_2855(g20627,g17433);
  IV  NOT_2856(I12837,g4222);
  IV  NOT_2857(g7892,g4801);
  IV  NOT_2858(g34934,g34918);
  IV  NOT_2859(g9558,g5841);
  IV  NOT_2860(g20379,g17821);
  IV  NOT_2861(g8057,g3068);
  IV  NOT_2862(g32564,g31376);
  IV  NOT_2863(I13995,g8744);
  IV  NOT_2864(g24379,g22550);
  IV  NOT_2865(g8457,g225);
  IV  NOT_2866(g8989,I12935);
  IV  NOT_2867(g19352,g15758);
  IV  NOT_2868(g22546,I21918);
  IV  NOT_2869(g23760,I22889);
  IV  NOT_2870(g20050,I20321);
  IV  NOT_2871(g23029,g20453);
  IV  NOT_2872(g6804,g490);
  IV  NOT_2873(g24112,g19935);
  IV  NOT_2874(g10367,g6870);
  IV  NOT_2875(g10394,g6994);
  IV  NOT_2876(I25028,g24484);
  IV  NOT_2877(g24050,g20841);
  IV  NOT_2878(g9901,g84);
  IV  NOT_2879(g34692,I32846);
  IV  NOT_2880(I22143,g20189);
  IV  NOT_2881(I21784,g19638);
  IV  NOT_2882(g23506,g21514);
  IV  NOT_2883(g23028,g20391);
  IV  NOT_2884(I18752,g6358);
  IV  NOT_2885(I28480,g28652);
  IV  NOT_2886(g31814,g29385);
  IV  NOT_2887(g32673,g31376);
  IV  NOT_2888(g32847,g30735);
  IV  NOT_2889(g20386,g15224);
  IV  NOT_2890(I21297,g18597);
  IV  NOT_2891(g8971,I12927);
  IV  NOT_2892(g22860,g20000);
  IV  NOT_2893(g24386,g22594);
  IV  NOT_2894(g20603,g17873);
  IV  NOT_2895(g9511,g5881);
  IV  NOT_2896(g27736,I26356);
  IV  NOT_2897(g7738,I12176);
  IV  NOT_2898(g31807,g29385);
  IV  NOT_2899(g8686,g2819);
  IV  NOT_2900(g13302,g12321);
  IV  NOT_2901(g20096,g16782);
  IV  NOT_2902(g24603,g23108);
  IV  NOT_2903(g33772,I31622);
  IV  NOT_2904(g7991,g4878);
  IV  NOT_2905(I23354,g23277);
  IV  NOT_2906(g24096,g19890);
  IV  NOT_2907(g29922,g28837);
  IV  NOT_2908(g34400,g34142);
  IV  NOT_2909(g7244,g4408);
  IV  NOT_2910(g12887,g10394);
  IV  NOT_2911(g10420,g9239);
  IV  NOT_2912(I17143,g14412);
  IV  NOT_2913(g22497,g19513);
  IV  NOT_2914(g25184,g22763);
  IV  NOT_2915(g32509,g31070);
  IV  NOT_2916(g31639,I29225);
  IV  NOT_2917(g10319,I13740);
  IV  NOT_2918(g17088,I18160);
  IV  NOT_2919(g32933,g31376);
  IV  NOT_2920(g30329,I28588);
  IV  NOT_2921(g9492,g2759);
  IV  NOT_2922(I21181,g17413);
  IV  NOT_2923(g16136,I17491);
  IV  NOT_2924(g7340,g4443);
  IV  NOT_2925(g20681,g15483);
  IV  NOT_2926(g9600,g3632);
  IV  NOT_2927(I23671,g23202);
  IV  NOT_2928(g32508,g30825);
  IV  NOT_2929(g9574,g6462);
  IV  NOT_2930(g31638,g29689);
  IV  NOT_2931(g9864,I13424);
  IV  NOT_2932(g32634,g30673);
  IV  NOT_2933(g32851,g31327);
  IV  NOT_2934(g32872,g31327);
  IV  NOT_2935(g33638,I31469);
  IV  NOT_2936(g35001,I33297);
  IV  NOT_2937(g30328,I28585);
  IV  NOT_2938(g7907,g3072);
  IV  NOT_2939(g11640,I14550);
  IV  NOT_2940(g11769,g8626);
  IV  NOT_2941(g34539,g34354);
  IV  NOT_2942(g9714,g4012);
  IV  NOT_2943(g12843,g10359);
  IV  NOT_2944(g17497,g14879);
  IV  NOT_2945(g22987,g20391);
  IV  NOT_2946(g34328,g34096);
  IV  NOT_2947(g10059,g6451);
  IV  NOT_2948(g23927,g19074);
  IV  NOT_2949(I18842,g13809);
  IV  NOT_2950(g24429,g22722);
  IV  NOT_2951(g19524,g15695);
  IV  NOT_2952(I29891,g31578);
  IV  NOT_2953(g7517,g962);
  IV  NOT_2954(g22658,I21969);
  IV  NOT_2955(g29953,g28907);
  IV  NOT_2956(g10540,g9392);
  IV  NOT_2957(g10058,g6497);
  IV  NOT_2958(g31841,g29385);
  IV  NOT_2959(g24428,g22722);
  IV  NOT_2960(I32096,g33641);
  IV  NOT_2961(g33391,g32384);
  IV  NOT_2962(g19477,g16431);
  IV  NOT_2963(g12869,g10376);
  IV  NOT_2964(g16164,I17507);
  IV  NOT_2965(g23649,g18833);
  IV  NOT_2966(g26683,g25514);
  IV  NOT_2967(g7876,g1495);
  IV  NOT_2968(g25692,I24839);
  IV  NOT_2969(g15614,g14914);
  IV  NOT_2970(g22339,g19801);
  IV  NOT_2971(g20765,g17748);
  IV  NOT_2972(g8938,g4899);
  IV  NOT_2973(I19235,g15078);
  IV  NOT_2974(I20495,g16283);
  IV  NOT_2975(g29800,g28363);
  IV  NOT_2976(g10203,g2393);
  IV  NOT_2977(g12868,g10377);
  IV  NOT_2978(g21903,I21480);
  IV  NOT_2979(g14203,g12381);
  IV  NOT_2980(g20549,g15277);
  IV  NOT_2981(g23648,g18833);
  IV  NOT_2982(g13881,I16181);
  IV  NOT_2983(I16090,g10430);
  IV  NOT_2984(g22338,g19801);
  IV  NOT_2985(g23491,g21514);
  IV  NOT_2986(I20816,g17088);
  IV  NOT_2987(g23903,g18997);
  IV  NOT_2988(I33252,g34974);
  IV  NOT_2989(I32681,g34429);
  IV  NOT_2990(g10044,g5357);
  IV  NOT_2991(g34241,I32222);
  IV  NOT_2992(g27709,I26337);
  IV  NOT_2993(g21604,g15938);
  IV  NOT_2994(I22580,g20982);
  IV  NOT_2995(I16651,g10542);
  IV  NOT_2996(g20548,g15426);
  IV  NOT_2997(g8519,g287);
  IV  NOT_2998(g8740,I12735);
  IV  NOT_2999(g31578,I29199);
  IV  NOT_3000(g25013,g23599);
  IV  NOT_3001(g31835,g29385);
  IV  NOT_3002(g32574,g31070);
  IV  NOT_3003(I20985,g16300);
  IV  NOT_3004(g24548,g22942);
  IV  NOT_3005(I31564,g33204);
  IV  NOT_3006(g17296,I18280);
  IV  NOT_3007(g25214,g22228);
  IV  NOT_3008(g27708,I26334);
  IV  NOT_3009(I12418,g55);
  IV  NOT_3010(g17644,g15002);
  IV  NOT_3011(g20504,g18008);
  IV  NOT_3012(g30100,g29131);
  IV  NOT_3013(g23563,g20682);
  IV  NOT_3014(g10377,g6940);
  IV  NOT_3015(g32912,g30735);
  IV  NOT_3016(g8606,g4653);
  IV  NOT_3017(I18865,g14314);
  IV  NOT_3018(I20954,g16228);
  IV  NOT_3019(g19748,g17015);
  IV  NOT_3020(g10120,g1902);
  IV  NOT_3021(g22197,g19074);
  IV  NOT_3022(g14377,g12201);
  IV  NOT_3023(I11753,g4492);
  IV  NOT_3024(g22855,g20391);
  IV  NOT_3025(g19276,g17367);
  IV  NOT_3026(g9889,g6128);
  IV  NOT_3027(g13027,I15647);
  IV  NOT_3028(g7110,g6682);
  IV  NOT_3029(I14660,g9746);
  IV  NOT_3030(g33442,g31937);
  IV  NOT_3031(g22870,g20887);
  IV  NOT_3032(g22527,g19546);
  IV  NOT_3033(I21860,g19638);
  IV  NOT_3034(g34683,I32827);
  IV  NOT_3035(g28127,g27102);
  IV  NOT_3036(g25538,g22594);
  IV  NOT_3037(g29216,I27564);
  IV  NOT_3038(I32690,g34432);
  IV  NOT_3039(g11249,g8405);
  IV  NOT_3040(I28838,g29372);
  IV  NOT_3041(I13031,g6747);
  IV  NOT_3042(g14738,I16821);
  IV  NOT_3043(g13249,g10590);
  IV  NOT_3044(g14562,g12036);
  IV  NOT_3045(g14645,I16755);
  IV  NOT_3046(I30861,g32383);
  IV  NOT_3047(g20129,g17328);
  IV  NOT_3048(g16606,g14110);
  IV  NOT_3049(g17197,I18233);
  IV  NOT_3050(g18880,g15656);
  IV  NOT_3051(g23767,g18997);
  IV  NOT_3052(g23794,g19147);
  IV  NOT_3053(g21395,g17873);
  IV  NOT_3054(g24129,g20857);
  IV  NOT_3055(g32592,g30673);
  IV  NOT_3056(g20057,g16349);
  IV  NOT_3057(g32756,g31021);
  IV  NOT_3058(g23395,I22502);
  IV  NOT_3059(g24057,g20841);
  IV  NOT_3060(g20128,g17533);
  IV  NOT_3061(I12167,g5176);
  IV  NOT_3062(g14290,I16460);
  IV  NOT_3063(g17870,I18842);
  IV  NOT_3064(g17411,g14454);
  IV  NOT_3065(g17527,g14741);
  IV  NOT_3066(g23899,g19277);
  IV  NOT_3067(g7002,g5160);
  IV  NOT_3068(g13003,I15609);
  IV  NOT_3069(g24128,g20720);
  IV  NOT_3070(g11204,I14271);
  IV  NOT_3071(I14550,g10072);
  IV  NOT_3072(g7824,g4169);
  IV  NOT_3073(g30991,I28925);
  IV  NOT_3074(g6996,g4955);
  IV  NOT_3075(g25241,g23651);
  IV  NOT_3076(g11779,g9602);
  IV  NOT_3077(I18270,g13191);
  IV  NOT_3078(g16750,g14454);
  IV  NOT_3079(g22867,g20391);
  IV  NOT_3080(g34991,I33273);
  IV  NOT_3081(g7236,g4608);
  IV  NOT_3082(g9285,g2715);
  IV  NOT_3083(g20626,g15483);
  IV  NOT_3084(g27774,I26381);
  IV  NOT_3085(I27401,g27051);
  IV  NOT_3086(I11843,g111);
  IV  NOT_3087(g23898,g19277);
  IV  NOT_3088(g9500,g5495);
  IV  NOT_3089(g20323,g17873);
  IV  NOT_3090(I21250,g16540);
  IV  NOT_3091(g29117,g27886);
  IV  NOT_3092(g24626,g23139);
  IV  NOT_3093(g33430,g32421);
  IV  NOT_3094(g23191,I22289);
  IV  NOT_3095(g20533,g17271);
  IV  NOT_3096(g10427,g10053);
  IV  NOT_3097(g12955,I15577);
  IV  NOT_3098(g32820,g31672);
  IV  NOT_3099(I18460,g5276);
  IV  NOT_3100(g8341,g3119);
  IV  NOT_3101(g10366,g6895);
  IV  NOT_3102(g24533,g22876);
  IV  NOT_3103(g25100,g22384);
  IV  NOT_3104(g12879,g10381);
  IV  NOT_3105(g22714,g20436);
  IV  NOT_3106(g11786,g7549);
  IV  NOT_3107(g14366,I16526);
  IV  NOT_3108(g17503,g14892);
  IV  NOT_3109(I14054,g10028);
  IV  NOT_3110(g9184,g6120);
  IV  NOT_3111(g23521,g21468);
  IV  NOT_3112(g28181,I26700);
  IV  NOT_3113(g25771,I24920);
  IV  NOT_3114(g20775,g18008);
  IV  NOT_3115(g18831,g15224);
  IV  NOT_3116(I15647,g12109);
  IV  NOT_3117(I23339,g23232);
  IV  NOT_3118(g32846,g31376);
  IV  NOT_3119(g9339,g2295);
  IV  NOT_3120(I19759,g17767);
  IV  NOT_3121(g19733,g16856);
  IV  NOT_3122(I24558,g23777);
  IV  NOT_3123(g12878,g10386);
  IV  NOT_3124(g26758,g25389);
  IV  NOT_3125(I27749,g28917);
  IV  NOT_3126(I20830,g17657);
  IV  NOT_3127(g12337,g9340);
  IV  NOT_3128(g32731,g31376);
  IV  NOT_3129(g31806,g29385);
  IV  NOT_3130(g22202,I21784);
  IV  NOT_3131(g33806,I31650);
  IV  NOT_3132(g9024,g4358);
  IV  NOT_3133(I12749,g4575);
  IV  NOT_3134(g11826,I14650);
  IV  NOT_3135(g17714,g14930);
  IV  NOT_3136(g12886,g10393);
  IV  NOT_3137(g22979,g20453);
  IV  NOT_3138(g20737,g15656);
  IV  NOT_3139(g22496,g19510);
  IV  NOT_3140(g10403,g7040);
  IV  NOT_3141(I21969,g21370);
  IV  NOT_3142(g23440,I22557);
  IV  NOT_3143(g13999,g11048);
  IV  NOT_3144(g7222,g4427);
  IV  NOT_3145(g27967,I26479);
  IV  NOT_3146(g27994,g26793);
  IV  NOT_3147(g33142,g32072);
  IV  NOT_3148(g19630,g16897);
  IV  NOT_3149(g9809,g6082);
  IV  NOT_3150(g20232,g16931);
  IV  NOT_3151(I14773,g9581);
  IV  NOT_3152(g29814,I28062);
  IV  NOT_3153(g17819,I18825);
  IV  NOT_3154(g17707,g14758);
  IV  NOT_3155(I33047,g34776);
  IV  NOT_3156(g30206,g28436);
  IV  NOT_3157(g7928,g4776);
  IV  NOT_3158(g26744,g25400);
  IV  NOT_3159(g12967,g11790);
  IV  NOT_3160(g23861,g19147);
  IV  NOT_3161(g23573,g20248);
  IV  NOT_3162(g32691,g30673);
  IV  NOT_3163(g18989,g16000);
  IV  NOT_3164(g8879,I12858);
  IV  NOT_3165(g8607,g37);
  IV  NOT_3166(g11233,g9664);
  IV  NOT_3167(I18875,g13782);
  IV  NOT_3168(g21247,g15171);
  IV  NOT_3169(g23247,g20924);
  IV  NOT_3170(g11182,I14241);
  IV  NOT_3171(I11708,g3703);
  IV  NOT_3172(g7064,g5990);
  IV  NOT_3173(g17818,I18822);
  IV  NOT_3174(g9672,g5390);
  IV  NOT_3175(I13708,g136);
  IV  NOT_3176(g20697,g17433);
  IV  NOT_3177(g14226,g11618);
  IV  NOT_3178(g9077,g504);
  IV  NOT_3179(g17496,g14683);
  IV  NOT_3180(I19345,g15083);
  IV  NOT_3181(g22986,g20330);
  IV  NOT_3182(g8659,g2815);
  IV  NOT_3183(g25882,g25026);
  IV  NOT_3184(g23926,g19074);
  IV  NOT_3185(g8358,I12541);
  IV  NOT_3186(g18988,g15979);
  IV  NOT_3187(I32775,g34512);
  IV  NOT_3188(g9477,I13149);
  IV  NOT_3189(g8506,g3782);
  IV  NOT_3190(I30766,g32363);
  IV  NOT_3191(g9523,g6419);
  IV  NOT_3192(g24995,g22763);
  IV  NOT_3193(g34759,I32935);
  IV  NOT_3194(g7785,g4621);
  IV  NOT_3195(g16522,g13889);
  IV  NOT_3196(g23612,I22745);
  IV  NOT_3197(g10572,g10233);
  IV  NOT_3198(I25534,g25448);
  IV  NOT_3199(I17964,g3661);
  IV  NOT_3200(g23388,g21070);
  IV  NOT_3201(I15932,g12381);
  IV  NOT_3202(g17590,I18523);
  IV  NOT_3203(g19476,g16326);
  IV  NOT_3204(g12919,I15536);
  IV  NOT_3205(I12808,g4322);
  IV  NOT_3206(g6799,g199);
  IV  NOT_3207(g26804,g25400);
  IV  NOT_3208(g20512,g18062);
  IV  NOT_3209(g34435,I32476);
  IV  NOT_3210(g23777,I22918);
  IV  NOT_3211(g23534,I22665);
  IV  NOT_3212(I26451,g26862);
  IV  NOT_3213(g13932,g11534);
  IV  NOT_3214(g32929,g31710);
  IV  NOT_3215(g8587,g3689);
  IV  NOT_3216(I14839,g9689);
  IV  NOT_3217(g23272,g20924);
  IV  NOT_3218(g11513,g7948);
  IV  NOT_3219(g19454,g16349);
  IV  NOT_3220(g7563,g6322);
  IV  NOT_3221(g17741,g12972);
  IV  NOT_3222(g12918,I15533);
  IV  NOT_3223(I18160,g14441);
  IV  NOT_3224(I15448,g10877);
  IV  NOT_3225(g17384,I18323);
  IV  NOT_3226(g32583,g30614);
  IV  NOT_3227(g32928,g31672);
  IV  NOT_3228(g19570,g16349);
  IV  NOT_3229(g19712,g17096);
  IV  NOT_3230(g6997,g4578);
  IV  NOT_3231(g22150,g21280);
  IV  NOT_3232(g11897,I14705);
  IV  NOT_3233(I22000,g20277);
  IV  NOT_3234(g10490,g9274);
  IV  NOT_3235(g9551,g3281);
  IV  NOT_3236(g9742,g6144);
  IV  NOT_3237(g9104,I12987);
  IV  NOT_3238(g23462,I22589);
  IV  NOT_3239(g9099,g3706);
  IV  NOT_3240(g34345,I32352);
  IV  NOT_3241(g9499,g5152);
  IV  NOT_3242(g11404,g7596);
  IV  NOT_3243(g15750,g13291);
  IV  NOT_3244(g34940,g34924);
  IV  NOT_3245(g13505,g10981);
  IV  NOT_3246(I15717,g6346);
  IV  NOT_3247(g16326,I17658);
  IV  NOT_3248(g18887,g15373);
  IV  NOT_3249(g20445,g15224);
  IV  NOT_3250(I31820,g33323);
  IV  NOT_3251(I12064,g617);
  IV  NOT_3252(g23032,I22211);
  IV  NOT_3253(g10376,g6923);
  IV  NOT_3254(g10385,I13805);
  IV  NOT_3255(g25206,g23613);
  IV  NOT_3256(g12598,g7004);
  IV  NOT_3257(g14376,g12126);
  IV  NOT_3258(g14385,I16541);
  IV  NOT_3259(g34848,I33070);
  IV  NOT_3260(g19074,I19772);
  IV  NOT_3261(g17735,g14807);
  IV  NOT_3262(g14297,g10869);
  IV  NOT_3263(g20499,g15483);
  IV  NOT_3264(g7394,g5637);
  IV  NOT_3265(g10980,g9051);
  IV  NOT_3266(g11026,g8434);
  IV  NOT_3267(I26785,g27013);
  IV  NOT_3268(g12086,g9654);
  IV  NOT_3269(g32787,g30937);
  IV  NOT_3270(g13026,g11018);
  IV  NOT_3271(g31863,I29447);
  IV  NOT_3272(I14619,g4185);
  IV  NOT_3273(g10354,g6811);
  IV  NOT_3274(I23315,g21685);
  IV  NOT_3275(I33152,g34900);
  IV  NOT_3276(g19567,g16164);
  IV  NOT_3277(g14095,g11326);
  IV  NOT_3278(g29014,g27742);
  IV  NOT_3279(g22526,g19801);
  IV  NOT_3280(I17569,g14564);
  IV  NOT_3281(g9754,g2020);
  IV  NOT_3282(g21061,I20929);
  IV  NOT_3283(g28126,g27122);
  IV  NOT_3284(g18528,I19348);
  IV  NOT_3285(g20498,g15348);
  IV  NOT_3286(g6802,g468);
  IV  NOT_3287(g8284,g5002);
  IV  NOT_3288(g23061,g20283);
  IV  NOT_3289(g8239,g1056);
  IV  NOT_3290(g28250,g27074);
  IV  NOT_3291(g10181,g2551);
  IV  NOT_3292(g25114,I24278);
  IV  NOT_3293(g7557,g1500);
  IV  NOT_3294(g8180,g262);
  IV  NOT_3295(I17747,g13298);
  IV  NOT_3296(g12322,I15162);
  IV  NOT_3297(g27977,g26105);
  IV  NOT_3298(g32743,g30937);
  IV  NOT_3299(g32827,g31672);
  IV  NOT_3300(g25082,g22342);
  IV  NOT_3301(g8591,g3763);
  IV  NOT_3302(g30332,I28597);
  IV  NOT_3303(g24056,g20014);
  IV  NOT_3304(g9613,g5062);
  IV  NOT_3305(g12901,g10404);
  IV  NOT_3306(g20611,g18008);
  IV  NOT_3307(g17526,I18469);
  IV  NOT_3308(g12977,I15590);
  IV  NOT_3309(g20080,g17328);
  IV  NOT_3310(g7471,g6012);
  IV  NOT_3311(g9044,g604);
  IV  NOT_3312(g20924,I20895);
  IV  NOT_3313(g19519,g16795);
  IV  NOT_3314(g24080,g21143);
  IV  NOT_3315(g19675,g16987);
  IV  NOT_3316(g9444,g5535);
  IV  NOT_3317(g9269,g5517);
  IV  NOT_3318(g22866,g20330);
  IV  NOT_3319(I17814,g3274);
  IV  NOT_3320(g32640,g31154);
  IV  NOT_3321(g20432,g17847);
  IV  NOT_3322(g32769,g31672);
  IV  NOT_3323(g23360,I22461);
  IV  NOT_3324(g29116,g27837);
  IV  NOT_3325(g19518,g16239);
  IV  NOT_3326(g8507,g3712);
  IV  NOT_3327(g9983,g4239);
  IV  NOT_3328(g12656,g7028);
  IV  NOT_3329(I15620,g12038);
  IV  NOT_3330(I17772,g14888);
  IV  NOT_3331(g25849,g24491);
  IV  NOT_3332(g9862,g5413);
  IV  NOT_3333(I27555,g28142);
  IV  NOT_3334(g23447,g21562);
  IV  NOT_3335(g32768,g30825);
  IV  NOT_3336(g32803,g31376);
  IV  NOT_3337(g25399,g22763);
  IV  NOT_3338(g12295,g7139);
  IV  NOT_3339(I23384,g23362);
  IV  NOT_3340(g10190,g6044);
  IV  NOT_3341(g29041,I27385);
  IV  NOT_3342(g13620,g10556);
  IV  NOT_3343(g12823,g9206);
  IV  NOT_3344(I17639,g13350);
  IV  NOT_3345(I27570,g28262);
  IV  NOT_3346(I15811,g11128);
  IV  NOT_3347(I21067,g15573);
  IV  NOT_3348(I18822,g13745);
  IV  NOT_3349(g16509,g13873);
  IV  NOT_3350(I32056,g33641);
  IV  NOT_3351(g11811,g9724);
  IV  NOT_3352(I12712,g59);
  IV  NOT_3353(g20145,g17533);
  IV  NOT_3354(g34833,I33047);
  IV  NOT_3355(g34049,g33678);
  IV  NOT_3356(I13010,g6749);
  IV  NOT_3357(g31821,g29385);
  IV  NOT_3358(g32881,g30673);
  IV  NOT_3359(I32988,g34755);
  IV  NOT_3360(g24031,g21193);
  IV  NOT_3361(I33020,g34781);
  IV  NOT_3362(g16508,I17704);
  IV  NOT_3363(I24455,g22541);
  IV  NOT_3364(g26605,g25293);
  IV  NOT_3365(g20650,g15348);
  IV  NOT_3366(g23629,g21514);
  IV  NOT_3367(g21451,I21162);
  IV  NOT_3368(g16872,I18060);
  IV  NOT_3369(I12907,g4322);
  IV  NOT_3370(g22923,I22124);
  IV  NOT_3371(I17416,g13806);
  IV  NOT_3372(g23472,g21062);
  IV  NOT_3373(g15483,I17128);
  IV  NOT_3374(g9534,g90);
  IV  NOT_3375(g9729,g5138);
  IV  NOT_3376(g9961,g6404);
  IV  NOT_3377(g7438,g5983);
  IV  NOT_3378(g25263,g22763);
  IV  NOT_3379(g29983,g28977);
  IV  NOT_3380(g20529,g15509);
  IV  NOT_3381(g22300,I21815);
  IV  NOT_3382(g26812,g25439);
  IV  NOT_3383(I21019,g17325);
  IV  NOT_3384(g27017,g25895);
  IV  NOT_3385(I27567,g28181);
  IV  NOT_3386(g15862,I17355);
  IV  NOT_3387(g8515,I12631);
  IV  NOT_3388(g34221,I32192);
  IV  NOT_3389(g8630,g4843);
  IV  NOT_3390(g21246,I20985);
  IV  NOT_3391(I27238,g27320);
  IV  NOT_3392(g23246,g20785);
  IV  NOT_3393(g20528,g15224);
  IV  NOT_3394(g20696,g17533);
  IV  NOT_3395(g25135,g22457);
  IV  NOT_3396(g20330,I20542);
  IV  NOT_3397(g9927,g5689);
  IV  NOT_3398(g32662,g30614);
  IV  NOT_3399(g8300,g1242);
  IV  NOT_3400(g32027,I29585);
  IV  NOT_3401(I32461,g34244);
  IV  NOT_3402(g19577,g16129);
  IV  NOT_3403(g17688,I18667);
  IV  NOT_3404(g9014,g3004);
  IV  NOT_3405(g20764,I20819);
  IV  NOT_3406(g10497,g10102);
  IV  NOT_3407(I25591,g25380);
  IV  NOT_3408(g32890,g30735);
  IV  NOT_3409(I33282,g34987);
  IV  NOT_3410(I27941,g28803);
  IV  NOT_3411(g9414,g2004);
  IV  NOT_3412(g7212,g6411);
  IV  NOT_3413(g19439,g15885);
  IV  NOT_3414(g9660,g3267);
  IV  NOT_3415(g9946,g6093);
  IV  NOT_3416(g20132,g16931);
  IV  NOT_3417(g24365,g22594);
  IV  NOT_3418(g20869,g15615);
  IV  NOT_3419(g13412,g11963);
  IV  NOT_3420(g23776,g21177);
  IV  NOT_3421(g34947,g34938);
  IV  NOT_3422(I12382,g47);
  IV  NOT_3423(g24132,g19890);
  IV  NOT_3424(g32482,g30614);
  IV  NOT_3425(g24869,I24041);
  IV  NOT_3426(g24960,g23716);
  IV  NOT_3427(g19438,g16249);
  IV  NOT_3428(I12519,g3447);
  IV  NOT_3429(g17157,g13350);
  IV  NOT_3430(I12176,g5523);
  IV  NOT_3431(g9903,g681);
  IV  NOT_3432(g13133,g11330);
  IV  NOT_3433(g32710,g30825);
  IV  NOT_3434(I12092,g790);
  IV  NOT_3435(g14700,g12512);
  IV  NOT_3436(g21355,g17821);
  IV  NOT_3437(g32552,g30825);
  IV  NOT_3438(g31834,g29385);
  IV  NOT_3439(g23355,g21070);
  IV  NOT_3440(g34812,I33024);
  IV  NOT_3441(g10658,I13979);
  IV  NOT_3442(g21370,g16323);
  IV  NOT_3443(g23859,g19074);
  IV  NOT_3444(g28819,I27271);
  IV  NOT_3445(g16311,g13273);
  IV  NOT_3446(g32779,g30937);
  IV  NOT_3447(I17442,g13638);
  IV  NOT_3448(g18878,g15426);
  IV  NOT_3449(g24161,I23327);
  IV  NOT_3450(g29130,g27907);
  IV  NOT_3451(I32696,g34434);
  IV  NOT_3452(I32843,g34499);
  IV  NOT_3453(g7993,I12333);
  IV  NOT_3454(g20709,g15426);
  IV  NOT_3455(g11011,g10274);
  IV  NOT_3456(g22854,g20330);
  IV  NOT_3457(g34951,g34941);
  IV  NOT_3458(g34972,I33232);
  IV  NOT_3459(g23858,g18997);
  IV  NOT_3460(g13011,I15623);
  IV  NOT_3461(I12935,g6753);
  IV  NOT_3462(g32778,g31021);
  IV  NOT_3463(g18886,g16000);
  IV  NOT_3464(I31803,g33176);
  IV  NOT_3465(g9036,g5084);
  IV  NOT_3466(I18313,g13350);
  IV  NOT_3467(g25221,g23653);
  IV  NOT_3468(I22275,g20127);
  IV  NOT_3469(g8440,g3431);
  IV  NOT_3470(g20708,g15426);
  IV  NOT_3471(g22763,I22046);
  IV  NOT_3472(g9679,g5475);
  IV  NOT_3473(g23172,I22275);
  IV  NOT_3474(g13716,I16090);
  IV  NOT_3475(I17615,g13251);
  IV  NOT_3476(g20087,g17249);
  IV  NOT_3477(g32786,g31021);
  IV  NOT_3478(g33726,I31581);
  IV  NOT_3479(I32960,g34653);
  IV  NOT_3480(g8123,g3808);
  IV  NOT_3481(g19566,g16136);
  IV  NOT_3482(g14338,I16502);
  IV  NOT_3483(g24087,g21143);
  IV  NOT_3484(I18276,g1075);
  IV  NOT_3485(I18285,g13638);
  IV  NOT_3486(g28590,g27724);
  IV  NOT_3487(g23844,g21308);
  IV  NOT_3488(g32647,g31154);
  IV  NOT_3489(g23394,I22499);
  IV  NOT_3490(I32868,g34579);
  IV  NOT_3491(g9831,g2269);
  IV  NOT_3492(g32945,g30937);
  IV  NOT_3493(g33436,I30962);
  IV  NOT_3494(g22660,g19140);
  IV  NOT_3495(g15509,I17136);
  IV  NOT_3496(I19012,g15060);
  IV  NOT_3497(g17763,g15011);
  IV  NOT_3498(g8666,g3703);
  IV  NOT_3499(g10060,g6541);
  IV  NOT_3500(I18900,g16767);
  IV  NOT_3501(g27976,g26703);
  IV  NOT_3502(g27985,g26131);
  IV  NOT_3503(I32161,g33791);
  IV  NOT_3504(g32826,g30825);
  IV  NOT_3505(g25273,g23978);
  IV  NOT_3506(g29863,g28410);
  IV  NOT_3507(g24043,g20982);
  IV  NOT_3508(g10197,g31);
  IV  NOT_3509(I21300,g18598);
  IV  NOT_3510(g22456,g19801);
  IV  NOT_3511(g12976,I15587);
  IV  NOT_3512(g15634,I17188);
  IV  NOT_3513(I23688,g23244);
  IV  NOT_3514(I23300,g21665);
  IV  NOT_3515(g14197,g12160);
  IV  NOT_3516(g32090,g31003);
  IV  NOT_3517(g9805,g5485);
  IV  NOT_3518(g9916,g3625);
  IV  NOT_3519(g19653,g16897);
  IV  NOT_3520(g33346,g32132);
  IV  NOT_3521(I18101,g13416);
  IV  NOT_3522(I32225,g34121);
  IV  NOT_3523(g10527,I13892);
  IV  NOT_3524(I12577,g1227);
  IV  NOT_3525(g10411,g7086);
  IV  NOT_3526(g23420,g21514);
  IV  NOT_3527(g9749,g1691);
  IV  NOT_3528(I18177,g13191);
  IV  NOT_3529(I18560,g5969);
  IV  NOT_3530(g32651,g31376);
  IV  NOT_3531(g18918,I19704);
  IV  NOT_3532(g32672,g31579);
  IV  NOT_3533(I19789,g17793);
  IV  NOT_3534(g24069,g19968);
  IV  NOT_3535(g22550,I21922);
  IV  NOT_3536(I33027,g34767);
  IV  NOT_3537(g26788,g25349);
  IV  NOT_3538(g26724,g25341);
  IV  NOT_3539(g20657,g17433);
  IV  NOT_3540(g20774,g18008);
  IV  NOT_3541(I26427,g26859);
  IV  NOT_3542(g8655,g2787);
  IV  NOT_3543(g23446,g21562);
  IV  NOT_3544(I16057,g10430);
  IV  NOT_3545(I28908,g30182);
  IV  NOT_3546(g19636,g16987);
  IV  NOT_3547(g23227,g20924);
  IV  NOT_3548(g30012,I28241);
  IV  NOT_3549(g19415,g15758);
  IV  NOT_3550(g24068,g19919);
  IV  NOT_3551(g24375,g22722);
  IV  NOT_3552(g21059,g15509);
  IV  NOT_3553(I33249,g34971);
  IV  NOT_3554(g7462,g2599);
  IV  NOT_3555(g23059,g20453);
  IV  NOT_3556(g31797,g29385);
  IV  NOT_3557(g6838,g1724);
  IV  NOT_3558(g13096,I15727);
  IV  NOT_3559(g33641,I31474);
  IV  NOT_3560(g32932,g31327);
  IV  NOT_3561(g33797,g33306);
  IV  NOT_3562(I31482,g33204);
  IV  NOT_3563(g19852,g17015);
  IV  NOT_3564(g22721,I22028);
  IV  NOT_3565(g10503,g8879);
  IV  NOT_3566(I16626,g11986);
  IV  NOT_3567(g21058,g15426);
  IV  NOT_3568(g6809,g341);
  IV  NOT_3569(g32513,g31376);
  IV  NOT_3570(I20864,g16960);
  IV  NOT_3571(g23058,g20453);
  IV  NOT_3572(g32449,I29977);
  IV  NOT_3573(g14503,g12256);
  IV  NOT_3574(g16691,g14160);
  IV  NOT_3575(I24022,g22182);
  IV  NOT_3576(g19963,g16326);
  IV  NOT_3577(g12842,g10355);
  IV  NOT_3578(g34473,g34426);
  IV  NOT_3579(I12083,g568);
  IV  NOT_3580(g17085,g14238);
  IV  NOT_3581(I31779,g33212);
  IV  NOT_3582(g24171,I23357);
  IV  NOT_3583(g32897,g30735);
  IV  NOT_3584(g32961,g31376);
  IV  NOT_3585(g23203,g20073);
  IV  NOT_3586(g8839,I12819);
  IV  NOT_3587(g34789,I32997);
  IV  NOT_3588(g7788,g4674);
  IV  NOT_3589(g11429,g7616);
  IV  NOT_3590(g17721,g12915);
  IV  NOT_3591(g29372,I27738);
  IV  NOT_3592(g10581,g9529);
  IV  NOT_3593(I16775,g12183);
  IV  NOT_3594(g13857,I16163);
  IV  NOT_3595(g32505,g31566);
  IV  NOT_3596(g20994,g15615);
  IV  NOT_3597(g9095,g3368);
  IV  NOT_3598(g32404,I29936);
  IV  NOT_3599(I14800,g10107);
  IV  NOT_3600(g33136,g32057);
  IV  NOT_3601(g9037,g164);
  IV  NOT_3602(g14714,g11405);
  IV  NOT_3603(g33635,g33436);
  IV  NOT_3604(g24994,g22432);
  IV  NOT_3605(g14315,I16479);
  IV  NOT_3606(g30325,I28576);
  IV  NOT_3607(g34788,I32994);
  IV  NOT_3608(g11793,I14633);
  IV  NOT_3609(g11428,g7615);
  IV  NOT_3610(g26682,g25309);
  IV  NOT_3611(g9653,g2441);
  IV  NOT_3612(g17431,I18376);
  IV  NOT_3613(g13793,I16120);
  IV  NOT_3614(g22341,g19801);
  IV  NOT_3615(g32717,g30735);
  IV  NOT_3616(g34325,g34092);
  IV  NOT_3617(I15765,g10823);
  IV  NOT_3618(I18009,g13680);
  IV  NOT_3619(g21281,g16286);
  IV  NOT_3620(g18977,g16100);
  IV  NOT_3621(I31786,g33197);
  IV  NOT_3622(I32970,g34716);
  IV  NOT_3623(g22156,g19147);
  IV  NOT_3624(g27830,g26802);
  IV  NOT_3625(g21902,I21477);
  IV  NOT_3626(g34920,I33152);
  IV  NOT_3627(g8172,g3873);
  IV  NOT_3628(g8278,g3096);
  IV  NOT_3629(g34434,I32473);
  IV  NOT_3630(g23902,g21468);
  IV  NOT_3631(g23301,g21037);
  IV  NOT_3632(g34358,I32364);
  IV  NOT_3633(g28917,I27314);
  IV  NOT_3634(g23377,g21070);
  IV  NOT_3635(I32878,g34501);
  IV  NOT_3636(g22180,g19210);
  IV  NOT_3637(g24425,g22722);
  IV  NOT_3638(g19554,g16861);
  IV  NOT_3639(g10111,g1858);
  IV  NOT_3640(g12830,g9995);
  IV  NOT_3641(g12893,g10391);
  IV  NOT_3642(I11816,g93);
  IV  NOT_3643(g16583,g14069);
  IV  NOT_3644(g7392,g4438);
  IV  NOT_3645(g20919,g15224);
  IV  NOT_3646(g15756,g13315);
  IV  NOT_3647(I25146,g24911);
  IV  NOT_3648(g34946,g34934);
  IV  NOT_3649(I25562,g25250);
  IV  NOT_3650(g19609,g16264);
  IV  NOT_3651(g8235,I12463);
  IV  NOT_3652(g8343,g3447);
  IV  NOT_3653(I18476,g14031);
  IV  NOT_3654(g34121,I32056);
  IV  NOT_3655(I14964,g10230);
  IV  NOT_3656(g19200,I19789);
  IV  NOT_3657(g21562,I21199);
  IV  NOT_3658(g9752,g1840);
  IV  NOT_3659(g12865,g10372);
  IV  NOT_3660(g20010,g17226);
  IV  NOT_3661(g8282,g3841);
  IV  NOT_3662(g20918,g15224);
  IV  NOT_3663(g23645,g20875);
  IV  NOT_3664(g8566,g3831);
  IV  NOT_3665(I18555,g5630);
  IV  NOT_3666(g24010,g21562);
  IV  NOT_3667(g9917,I13473);
  IV  NOT_3668(I32967,g34648);
  IV  NOT_3669(I32994,g34739);
  IV  NOT_3670(g10741,g8411);
  IV  NOT_3671(I21480,g18696);
  IV  NOT_3672(g7854,g1152);
  IV  NOT_3673(g13504,g11303);
  IV  NOT_3674(g25541,g22763);
  IV  NOT_3675(g20545,g15373);
  IV  NOT_3676(g20079,g17328);
  IV  NOT_3677(g20444,g15373);
  IV  NOT_3678(g21290,I21029);
  IV  NOT_3679(g32723,g31327);
  IV  NOT_3680(I31672,g33149);
  IV  NOT_3681(g10384,I13802);
  IV  NOT_3682(g8134,I12415);
  IV  NOT_3683(g23290,g20924);
  IV  NOT_3684(I33182,g34910);
  IV  NOT_3685(I13374,g6490);
  IV  NOT_3686(g8334,g3034);
  IV  NOT_3687(g24079,g20998);
  IV  NOT_3688(g21698,g18562);
  IV  NOT_3689(g14384,I16538);
  IV  NOT_3690(g22667,g21156);
  IV  NOT_3691(g34682,I32824);
  IV  NOT_3692(g29209,I27543);
  IV  NOT_3693(g20599,g18065);
  IV  NOT_3694(g6926,g3853);
  IV  NOT_3695(I16512,g12811);
  IV  NOT_3696(g23698,g21611);
  IV  NOT_3697(I12415,g48);
  IV  NOT_3698(g11317,I14346);
  IV  NOT_3699(g20078,g16846);
  IV  NOT_3700(I12333,g45);
  IV  NOT_3701(g32433,I29961);
  IV  NOT_3702(g19745,g16877);
  IV  NOT_3703(g24078,g20857);
  IV  NOT_3704(g6754,I11617);
  IV  NOT_3705(g12705,g7051);
  IV  NOT_3706(g20598,g17929);
  IV  NOT_3707(g32620,g30673);
  IV  NOT_3708(I28579,g29474);
  IV  NOT_3709(g20086,I20355);
  IV  NOT_3710(g19799,g17062);
  IV  NOT_3711(g25325,g22228);
  IV  NOT_3712(I32458,g34243);
  IV  NOT_3713(g11129,g7994);
  IV  NOT_3714(I25366,g24477);
  IV  NOT_3715(g8804,g4035);
  IV  NOT_3716(g10150,g1700);
  IV  NOT_3717(g24086,g20998);
  IV  NOT_3718(g16743,g13986);
  IV  NOT_3719(g21427,g17367);
  IV  NOT_3720(g15731,g13326);
  IV  NOT_3721(g9364,g5041);
  IV  NOT_3722(g10877,I14079);
  IV  NOT_3723(g23427,I22542);
  IV  NOT_3724(g25535,g22763);
  IV  NOT_3725(g32811,g30735);
  IV  NOT_3726(I12963,g640);
  IV  NOT_3727(g14150,g12381);
  IV  NOT_3728(g21366,I21100);
  IV  NOT_3729(g32646,g31070);
  IV  NOT_3730(g8792,I12790);
  IV  NOT_3731(g7219,g4405);
  IV  NOT_3732(g19798,g17200);
  IV  NOT_3733(I28014,g28158);
  IV  NOT_3734(g11128,g7993);
  IV  NOT_3735(g7640,I12128);
  IV  NOT_3736(I18238,g13144);
  IV  NOT_3737(g10019,g6479);
  IV  NOT_3738(g28157,I26670);
  IV  NOT_3739(I15626,g12041);
  IV  NOT_3740(g22210,I21792);
  IV  NOT_3741(g20322,g17873);
  IV  NOT_3742(g32971,g31672);
  IV  NOT_3743(g7431,g2555);
  IV  NOT_3744(I32079,g33937);
  IV  NOT_3745(g7252,g1592);
  IV  NOT_3746(g16640,I17834);
  IV  NOT_3747(g29913,g28840);
  IV  NOT_3748(g34760,I32938);
  IV  NOT_3749(g7812,I12214);
  IV  NOT_3750(g16769,g13530);
  IV  NOT_3751(g20159,g17533);
  IV  NOT_3752(g34134,I32079);
  IV  NOT_3753(g25121,g22432);
  IV  NOT_3754(g20901,I20867);
  IV  NOT_3755(g13626,g11273);
  IV  NOT_3756(g20532,g15277);
  IV  NOT_3757(g17487,I18414);
  IV  NOT_3758(I27576,g28173);
  IV  NOT_3759(I15533,g11867);
  IV  NOT_3760(g24159,I23321);
  IV  NOT_3761(g13323,g11048);
  IV  NOT_3762(g24125,g19890);
  IV  NOT_3763(g6983,g4698);
  IV  NOT_3764(I18382,g13350);
  IV  NOT_3765(g21661,I21222);
  IV  NOT_3766(g17502,g14697);
  IV  NOT_3767(g16768,g13223);
  IV  NOT_3768(I19927,g17408);
  IV  NOT_3769(g20158,g16971);
  IV  NOT_3770(g8113,g3466);
  IV  NOT_3771(g12938,I15556);
  IV  NOT_3772(I16498,g10430);
  IV  NOT_3773(g23403,I22512);
  IV  NOT_3774(g23547,g21611);
  IV  NOT_3775(g23895,g19147);
  IV  NOT_3776(I13424,g5689);
  IV  NOT_3777(g24158,I23318);
  IV  NOT_3778(g33750,I31607);
  IV  NOT_3779(I18092,g3668);
  IV  NOT_3780(g7405,g1936);
  IV  NOT_3781(g13298,I15862);
  IV  NOT_3782(g19732,g17096);
  IV  NOT_3783(I22264,g20100);
  IV  NOT_3784(I30980,g32132);
  IV  NOT_3785(I24008,g22182);
  IV  NOT_3786(g29905,g28783);
  IV  NOT_3787(g20561,g17873);
  IV  NOT_3788(g20656,g17249);
  IV  NOT_3789(g9553,I13202);
  IV  NOT_3790(I18518,g13835);
  IV  NOT_3791(I18154,g13177);
  IV  NOT_3792(g23226,g20924);
  IV  NOT_3793(g7765,g4165);
  IV  NOT_3794(g20680,g15348);
  IV  NOT_3795(g26648,g25115);
  IV  NOT_3796(g20144,g17533);
  IV  NOT_3797(g10402,g7023);
  IV  NOT_3798(g23715,g20764);
  IV  NOT_3799(g23481,I22604);
  IV  NOT_3800(g32850,g30937);
  IV  NOT_3801(g31796,g29385);
  IV  NOT_3802(g19761,g17015);
  IV  NOT_3803(I12608,g1582);
  IV  NOT_3804(g12875,I15494);
  IV  NOT_3805(I21734,g19268);
  IV  NOT_3806(g6961,I11734);
  IV  NOT_3807(g8567,g4082);
  IV  NOT_3808(I21930,g21297);
  IV  NOT_3809(g34927,I33173);
  IV  NOT_3810(g7733,g4093);
  IV  NOT_3811(I22422,g19330);
  IV  NOT_3812(I15697,g6000);
  IV  NOT_3813(I17873,g15017);
  IV  NOT_3814(g31840,g29385);
  IV  NOT_3815(I32158,g33791);
  IV  NOT_3816(g12218,I15073);
  IV  NOT_3817(g32896,g31376);
  IV  NOT_3818(g12837,g10354);
  IV  NOT_3819(g23127,g21163);
  IV  NOT_3820(g6927,g3845);
  IV  NOT_3821(I21838,g19263);
  IV  NOT_3822(g25134,g22417);
  IV  NOT_3823(g10001,g6105);
  IV  NOT_3824(g22975,g20391);
  IV  NOT_3825(g13856,I16160);
  IV  NOT_3826(I23694,g23252);
  IV  NOT_3827(I29248,g29491);
  IV  NOT_3828(g9888,g5831);
  IV  NOT_3829(g10077,g1724);
  IV  NOT_3830(g13995,g11261);
  IV  NOT_3831(I33149,g34900);
  IV  NOT_3832(g8593,g3759);
  IV  NOT_3833(g29153,g27937);
  IV  NOT_3834(g24966,g22763);
  IV  NOT_3835(g7073,g6191);
  IV  NOT_3836(I12799,g59);
  IV  NOT_3837(g20631,g15171);
  IV  NOT_3838(g17815,g14348);
  IV  NOT_3839(g10597,g10233);
  IV  NOT_3840(g23490,g21514);
  IV  NOT_3841(g25506,g22228);
  IV  NOT_3842(g9429,g3723);
  IV  NOT_3843(I13705,g63);
  IV  NOT_3844(I29204,g29505);
  IV  NOT_3845(g32716,g31376);
  IV  NOT_3846(g7473,g6697);
  IV  NOT_3847(g16249,I17590);
  IV  NOT_3848(g18976,g16100);
  IV  NOT_3849(g14597,I16713);
  IV  NOT_3850(g19539,g16129);
  IV  NOT_3851(g6946,I11721);
  IV  NOT_3852(g24017,g18833);
  IV  NOT_3853(g11512,g7634);
  IV  NOT_3854(g34648,I32752);
  IV  NOT_3855(g24364,g22722);
  IV  NOT_3856(g17677,g14882);
  IV  NOT_3857(g34491,I32550);
  IV  NOT_3858(I22542,g19773);
  IV  NOT_3859(g16482,g13464);
  IV  NOT_3860(I17834,g14977);
  IV  NOT_3861(g31522,I29185);
  IV  NOT_3862(g32582,g31170);
  IV  NOT_3863(g7980,g3161);
  IV  NOT_3864(g21297,I21042);
  IV  NOT_3865(g18954,g17427);
  IV  NOT_3866(g23376,g21070);
  IV  NOT_3867(g23385,I22488);
  IV  NOT_3868(I25095,g25265);
  IV  NOT_3869(g19538,g16100);
  IV  NOT_3870(g6903,g3502);
  IV  NOT_3871(g7069,g6137);
  IV  NOT_3872(g9281,I13057);
  IV  NOT_3873(I12805,g4098);
  IV  NOT_3874(g26990,g26105);
  IV  NOT_3875(g34755,I32929);
  IV  NOT_3876(g23889,g20682);
  IV  NOT_3877(I13124,g2729);
  IV  NOT_3878(I18728,g6012);
  IV  NOT_3879(I21210,g17526);
  IV  NOT_3880(g23354,g20453);
  IV  NOT_3881(I14579,g8792);
  IV  NOT_3882(g22169,g19147);
  IV  NOT_3883(I26700,g27956);
  IV  NOT_3884(g34770,I32956);
  IV  NOT_3885(g12470,I15284);
  IV  NOT_3886(g7540,I12026);
  IV  NOT_3887(g8160,g3423);
  IV  NOT_3888(g22884,g20453);
  IV  NOT_3889(g34981,g34973);
  IV  NOT_3890(g23888,g18997);
  IV  NOT_3891(g23824,g21271);
  IV  NOT_3892(I15831,g10416);
  IV  NOT_3893(g32627,g30673);
  IV  NOT_3894(g28307,g27306);
  IV  NOT_3895(g32959,g30937);
  IV  NOT_3896(g32925,g31327);
  IV  NOT_3897(g21181,g15426);
  IV  NOT_3898(g22168,g19147);
  IV  NOT_3899(g10102,g6727);
  IV  NOT_3900(g10157,g2036);
  IV  NOT_3901(g31862,I29444);
  IV  NOT_3902(g32958,g31710);
  IV  NOT_3903(I15316,g10087);
  IV  NOT_3904(I19719,g17431);
  IV  NOT_3905(g8450,g3821);
  IV  NOT_3906(g24023,g21127);
  IV  NOT_3907(g26718,g25168);
  IV  NOT_3908(I32364,g34208);
  IV  NOT_3909(g17791,g14950);
  IV  NOT_3910(g20571,g15277);
  IV  NOT_3911(g9684,g6191);
  IV  NOT_3912(g11316,g8967);
  IV  NOT_3913(g9745,g6537);
  IV  NOT_3914(g12075,I14935);
  IV  NOT_3915(I17436,g13416);
  IV  NOT_3916(g28431,I26925);
  IV  NOT_3917(g9639,g1752);
  IV  NOT_3918(I18906,g16963);
  IV  NOT_3919(g9338,g1870);
  IV  NOT_3920(g24571,g22942);
  IV  NOT_3921(g10231,g2661);
  IV  NOT_3922(I18083,g13394);
  IV  NOT_3923(g9963,g7);
  IV  NOT_3924(I26296,g26820);
  IV  NOT_3925(g33326,g32318);
  IV  NOT_3926(g17410,g12955);
  IV  NOT_3927(I12761,g4188);
  IV  NOT_3928(g11498,I14475);
  IV  NOT_3929(g34767,I32947);
  IV  NOT_3930(g14231,g12246);
  IV  NOT_3931(g26832,g24850);
  IV  NOT_3932(g34845,g34773);
  IV  NOT_3933(g32603,g31070);
  IV  NOT_3934(g6831,g1413);
  IV  NOT_3935(I22464,g21222);
  IV  NOT_3936(g23931,g20875);
  IV  NOT_3937(g32742,g31021);
  IV  NOT_3938(I29233,g30295);
  IV  NOT_3939(g9309,g5462);
  IV  NOT_3940(I23306,g21673);
  IV  NOT_3941(g30990,g29676);
  IV  NOT_3942(I18304,g14790);
  IV  NOT_3943(g19771,g17096);
  IV  NOT_3944(g25240,g23650);
  IV  NOT_3945(g32944,g31021);
  IV  NOT_3946(I29182,g30012);
  IV  NOT_3947(g29474,I27758);
  IV  NOT_3948(g34990,I33270);
  IV  NOT_3949(g11989,I14839);
  IV  NOT_3950(I25190,g25423);
  IV  NOT_3951(g16826,I18034);
  IV  NOT_3952(g17479,g14855);
  IV  NOT_3953(g21426,g15277);
  IV  NOT_3954(g8179,g4999);
  IV  NOT_3955(g12037,I14893);
  IV  NOT_3956(g20495,g17926);
  IV  NOT_3957(g23426,I22539);
  IV  NOT_3958(g25903,I25005);
  IV  NOT_3959(g27984,g26737);
  IV  NOT_3960(I13875,g1233);
  IV  NOT_3961(g33702,I31545);
  IV  NOT_3962(g9808,g5827);
  IV  NOT_3963(g19683,g16931);
  IV  NOT_3964(g23190,I22286);
  IV  NOT_3965(I16709,g10430);
  IV  NOT_3966(g11988,I14836);
  IV  NOT_3967(I21815,g21308);
  IV  NOT_3968(g17478,g14996);
  IV  NOT_3969(g28156,I26667);
  IV  NOT_3970(I12013,g590);
  IV  NOT_3971(g17015,I18143);
  IV  NOT_3972(g32681,g30735);
  IV  NOT_3973(I32309,g34210);
  IV  NOT_3974(I12214,g6561);
  IV  NOT_3975(g16182,g13846);
  IV  NOT_3976(g16651,g14005);
  IV  NOT_3977(I22153,g20014);
  IV  NOT_3978(g23520,g21468);
  IV  NOT_3979(g27155,g26131);
  IV  NOT_3980(g9759,g2265);
  IV  NOT_3981(g18830,g18008);
  IV  NOT_3982(I16471,g12367);
  IV  NOT_3983(g17486,I18411);
  IV  NOT_3984(g7898,g4991);
  IV  NOT_3985(g25563,g22594);
  IV  NOT_3986(g32802,g31327);
  IV  NOT_3987(g32857,g30937);
  IV  NOT_3988(g22223,g19210);
  IV  NOT_3989(g13271,I15834);
  IV  NOT_3990(g34718,I32884);
  IV  NOT_3991(g24985,g23586);
  IV  NOT_3992(g34521,g34270);
  IV  NOT_3993(g32730,g31327);
  IV  NOT_3994(g23546,g21611);
  IV  NOT_3995(I24215,g22360);
  IV  NOT_3996(g32793,g31021);
  IV  NOT_3997(I18653,g5681);
  IV  NOT_3998(g20374,g18065);
  IV  NOT_3999(g23211,g21308);
  IV  NOT_4000(I30644,g32024);
  IV  NOT_4001(g19882,g16540);
  IV  NOT_4002(g19414,g16349);
  IV  NOT_4003(g26701,g25341);
  IV  NOT_4004(g7245,I11896);
  IV  NOT_4005(g17580,I18509);
  IV  NOT_4006(g11753,g8587);
  IV  NOT_4007(I29961,g30984);
  IV  NOT_4008(I12538,g58);
  IV  NOT_4009(g26777,g25439);
  IV  NOT_4010(g20643,g15962);
  IV  NOT_4011(I18138,g14277);
  IV  NOT_4012(g9049,g640);
  IV  NOT_4013(g23088,I22240);
  IV  NOT_4014(g31847,g29385);
  IV  NOT_4015(g32765,g31327);
  IV  NOT_4016(g19407,g16268);
  IV  NOT_4017(g9449,g5770);
  IV  NOT_4018(g16449,I17679);
  IV  NOT_4019(g11031,g8609);
  IV  NOT_4020(g22922,g20330);
  IV  NOT_4021(g23860,g19074);
  IV  NOT_4022(I15650,g12110);
  IV  NOT_4023(g32690,g31070);
  IV  NOT_4024(g9575,g6509);
  IV  NOT_4025(g32549,g31554);
  IV  NOT_4026(I15736,g12322);
  IV  NOT_4027(I14684,g7717);
  IV  NOT_4028(I18333,g1083);
  IV  NOT_4029(g22179,g19210);
  IV  NOT_4030(I29717,g30931);
  IV  NOT_4031(g25262,g22763);
  IV  NOT_4032(I11617,g1);
  IV  NOT_4033(g11736,g8165);
  IV  NOT_4034(g20669,g15426);
  IV  NOT_4035(I17136,g14398);
  IV  NOT_4036(g16897,I18083);
  IV  NOT_4037(I26503,g26811);
  IV  NOT_4038(g34573,I32645);
  IV  NOT_4039(g7344,g5659);
  IV  NOT_4040(g25899,g24997);
  IV  NOT_4041(g13736,g11313);
  IV  NOT_4042(g32548,g30673);
  IV  NOT_4043(I18852,g13716);
  IV  NOT_4044(I32687,g34431);
  IV  NOT_4045(g34247,I32240);
  IV  NOT_4046(I32976,g34699);
  IV  NOT_4047(I32985,g34736);
  IV  NOT_4048(g22178,g19147);
  IV  NOT_4049(g9498,g5101);
  IV  NOT_4050(g6873,g3151);
  IV  NOT_4051(g20668,g15426);
  IV  NOT_4052(g34926,I33170);
  IV  NOT_4053(g32504,g30673);
  IV  NOT_4054(g31851,g29385);
  IV  NOT_4055(I15843,g11181);
  IV  NOT_4056(I32752,g34510);
  IV  NOT_4057(g9833,g2449);
  IV  NOT_4058(g10287,I13715);
  IV  NOT_4059(g7259,g4375);
  IV  NOT_4060(g21659,g17727);
  IV  NOT_4061(I33050,g34777);
  IV  NOT_4062(g14314,I16476);
  IV  NOT_4063(g16717,g13951);
  IV  NOT_4064(g17531,I18476);
  IV  NOT_4065(g12836,g10351);
  IV  NOT_4066(g20195,g16931);
  IV  NOT_4067(I26581,g26942);
  IV  NOT_4068(g8997,g577);
  IV  NOT_4069(g23987,g19277);
  IV  NOT_4070(g10085,g1768);
  IV  NOT_4071(g8541,g3498);
  IV  NOT_4072(g23250,g21070);
  IV  NOT_4073(g24489,I23694);
  IV  NOT_4074(I23363,g23385);
  IV  NOT_4075(g14307,I16468);
  IV  NOT_4076(I27235,g27320);
  IV  NOT_4077(g17178,I18214);
  IV  NOT_4078(g6869,I11691);
  IV  NOT_4079(g34777,I32973);
  IV  NOT_4080(g12477,I15295);
  IV  NOT_4081(g20525,g17955);
  IV  NOT_4082(I15869,g11234);
  IV  NOT_4083(g18939,g16077);
  IV  NOT_4084(g8132,I12411);
  IV  NOT_4085(g28443,I26936);
  IV  NOT_4086(g34272,g34229);
  IV  NOT_4087(g24525,g22670);
  IV  NOT_4088(g24424,g22722);
  IV  NOT_4089(I11623,g28);
  IV  NOT_4090(g13132,g10632);
  IV  NOT_4091(g17685,I18662);
  IV  NOT_4092(g17676,g12941);
  IV  NOT_4093(g13869,g10831);
  IV  NOT_4094(g20558,I20650);
  IV  NOT_4095(g8680,g686);
  IV  NOT_4096(g22936,g20283);
  IV  NOT_4097(I13623,g4294);
  IV  NOT_4098(I21486,g18727);
  IV  NOT_4099(g17953,I18861);
  IV  NOT_4100(I22327,g19367);
  IV  NOT_4101(g23339,g21070);
  IV  NOT_4102(g8353,I12530);
  IV  NOT_4103(g18938,g16053);
  IV  NOT_4104(g23943,g19147);
  IV  NOT_4105(g18093,I18885);
  IV  NOT_4106(I13037,g4304);
  IV  NOT_4107(I29149,g29384);
  IV  NOT_4108(g14431,g12208);
  IV  NOT_4109(g31213,I29013);
  IV  NOT_4110(g11868,g9185);
  IV  NOT_4111(g12864,g10373);
  IV  NOT_4112(g13868,g11493);
  IV  NOT_4113(g6917,g3684);
  IV  NOT_4114(g8744,g691);
  IV  NOT_4115(g23338,g20453);
  IV  NOT_4116(g18065,I18875);
  IV  NOT_4117(g24893,I24060);
  IV  NOT_4118(g12749,g7074);
  IV  NOT_4119(g19435,g16449);
  IV  NOT_4120(g9162,g622);
  IV  NOT_4121(g9019,I12950);
  IV  NOT_4122(g17417,g14804);
  IV  NOT_4123(I18609,g5976);
  IV  NOT_4124(g7886,g1442);
  IV  NOT_4125(g20544,g15171);
  IV  NOT_4126(g23969,g19277);
  IV  NOT_4127(g32626,g30614);
  IV  NOT_4128(g28039,g26365);
  IV  NOT_4129(I32195,g33628);
  IV  NOT_4130(I13352,g4146);
  IV  NOT_4131(g11709,I14584);
  IV  NOT_4132(g30997,g29702);
  IV  NOT_4133(g10156,g2675);
  IV  NOT_4134(g20713,g15277);
  IV  NOT_4135(g21060,g15509);
  IV  NOT_4136(g34997,I33291);
  IV  NOT_4137(I12991,g6752);
  IV  NOT_4138(g23060,g19908);
  IV  NOT_4139(g23968,g18833);
  IV  NOT_4140(g18875,g15171);
  IV  NOT_4141(g32533,g30614);
  IV  NOT_4142(g8558,g3787);
  IV  NOT_4143(g28038,g26365);
  IV  NOT_4144(I32525,g34285);
  IV  NOT_4145(g13259,I15824);
  IV  NOT_4146(g33912,I31770);
  IV  NOT_4147(g19744,g15885);
  IV  NOT_4148(g16620,I17808);
  IV  NOT_4149(g7314,g1740);
  IV  NOT_4150(g10180,g2259);
  IV  NOT_4151(I14006,g9104);
  IV  NOT_4152(I17108,g13782);
  IV  NOT_4153(I14475,g10175);
  IV  NOT_4154(g11471,g7626);
  IV  NOT_4155(g19345,g17591);
  IV  NOT_4156(g25099,g22369);
  IV  NOT_4157(g13087,g12012);
  IV  NOT_4158(g32775,g30825);
  IV  NOT_4159(g25388,g22763);
  IV  NOT_4160(g25324,g22228);
  IV  NOT_4161(I14727,g7753);
  IV  NOT_4162(g13258,I15821);
  IV  NOT_4163(g12900,g10406);
  IV  NOT_4164(g19399,g16489);
  IV  NOT_4165(g20610,g18008);
  IV  NOT_4166(g7870,g1193);
  IV  NOT_4167(g21411,g15426);
  IV  NOT_4168(g17762,g13000);
  IV  NOT_4169(g20705,I20793);
  IV  NOT_4170(g34766,g34703);
  IV  NOT_4171(g23870,g21293);
  IV  NOT_4172(I16010,g11148);
  IV  NOT_4173(g23411,g20734);
  IV  NOT_4174(g23527,g21611);
  IV  NOT_4175(g28187,I26710);
  IV  NOT_4176(I14222,g8286);
  IV  NOT_4177(I21922,g21335);
  IV  NOT_4178(g25534,g22763);
  IV  NOT_4179(g15932,I17395);
  IV  NOT_4180(g25098,g22369);
  IV  NOT_4181(g10335,g4483);
  IV  NOT_4182(I23321,g21693);
  IV  NOT_4183(g7650,g4064);
  IV  NOT_4184(g27101,g26770);
  IV  NOT_4185(g25272,g23715);
  IV  NOT_4186(g29862,g28406);
  IV  NOT_4187(g24042,g20014);
  IV  NOT_4188(g33072,g31945);
  IV  NOT_4189(g20189,I20447);
  IV  NOT_4190(g19398,g16489);
  IV  NOT_4191(g20679,g15634);
  IV  NOT_4192(I29368,g30321);
  IV  NOT_4193(g17423,I18360);
  IV  NOT_4194(g16971,I18131);
  IV  NOT_4195(g11043,g8561);
  IV  NOT_4196(g12036,g9245);
  IV  NOT_4197(g9086,g847);
  IV  NOT_4198(g32737,g31327);
  IV  NOT_4199(I18813,g5673);
  IV  NOT_4200(g17216,g14454);
  IV  NOT_4201(g20270,g15277);
  IV  NOT_4202(g9728,g5109);
  IV  NOT_4203(g19652,g16897);
  IV  NOT_4204(I30986,g32437);
  IV  NOT_4205(I17750,g14383);
  IV  NOT_4206(g22543,g19801);
  IV  NOT_4207(g17587,I18518);
  IV  NOT_4208(g9730,g5436);
  IV  NOT_4209(I31504,g33164);
  IV  NOT_4210(g24124,g21209);
  IV  NOT_4211(g8092,g1589);
  IV  NOT_4212(g14694,I16795);
  IV  NOT_4213(g29948,g28853);
  IV  NOT_4214(g8492,g3396);
  IV  NOT_4215(g9185,I13007);
  IV  NOT_4216(g23503,g21468);
  IV  NOT_4217(g23894,g19074);
  IV  NOT_4218(g19263,I19799);
  IV  NOT_4219(g32697,g31070);
  IV  NOT_4220(g27064,I25786);
  IV  NOT_4221(I18674,g13101);
  IV  NOT_4222(g25032,g23639);
  IV  NOT_4223(g20383,g15373);
  IV  NOT_4224(g32856,g31021);
  IV  NOT_4225(I28913,g30322);
  IV  NOT_4226(g11810,g9664);
  IV  NOT_4227(g25140,g22228);
  IV  NOT_4228(g9070,g5428);
  IV  NOT_4229(g8714,g4859);
  IV  NOT_4230(g7594,I12064);
  IV  NOT_4231(g31820,g29385);
  IV  NOT_4232(g10487,g10233);
  IV  NOT_4233(g32880,g30614);
  IV  NOT_4234(g13068,I15697);
  IV  NOT_4235(g25997,I25095);
  IV  NOT_4236(g7972,g1046);
  IV  NOT_4237(g24030,g21127);
  IV  NOT_4238(g20267,g17955);
  IV  NOT_4239(g24093,g20998);
  IV  NOT_4240(g10502,g8876);
  IV  NOT_4241(g26776,g25498);
  IV  NOT_4242(g23714,g20751);
  IV  NOT_4243(I27758,g28119);
  IV  NOT_4244(g23450,I22571);
  IV  NOT_4245(I29228,g30314);
  IV  NOT_4246(g32512,g31566);
  IV  NOT_4247(g7806,g4681);
  IV  NOT_4248(I15878,g11249);
  IV  NOT_4249(g20065,g16846);
  IV  NOT_4250(g31846,g29385);
  IV  NOT_4251(g7943,g1395);
  IV  NOT_4252(g24065,g20982);
  IV  NOT_4253(g11878,I14690);
  IV  NOT_4254(g19361,I19843);
  IV  NOT_4255(I20609,g16539);
  IV  NOT_4256(I12758,g4093);
  IV  NOT_4257(g23819,g19147);
  IV  NOT_4258(g12874,g10383);
  IV  NOT_4259(g26754,g25300);
  IV  NOT_4260(g34472,I32525);
  IV  NOT_4261(g25766,g24439);
  IV  NOT_4262(g28479,g27654);
  IV  NOT_4263(I32678,g34428);
  IV  NOT_4264(g23202,I22302);
  IV  NOT_4265(g14443,I16596);
  IV  NOT_4266(g23257,g20924);
  IV  NOT_4267(g26859,I25591);
  IV  NOT_4268(g27009,g25911);
  IV  NOT_4269(g26825,I25541);
  IV  NOT_4270(g21055,g15224);
  IV  NOT_4271(g23496,g20248);
  IV  NOT_4272(g7322,g1862);
  IV  NOT_4273(g16228,I17569);
  IV  NOT_4274(g20219,I20495);
  IV  NOT_4275(g23055,g20887);
  IV  NOT_4276(g6990,g4742);
  IV  NOT_4277(g17242,g14454);
  IV  NOT_4278(g34246,I32237);
  IV  NOT_4279(g10278,g4628);
  IV  NOT_4280(g33413,g31971);
  IV  NOT_4281(g29847,g28395);
  IV  NOT_4282(I29582,g30591);
  IV  NOT_4283(g23111,g20391);
  IV  NOT_4284(g12009,I14862);
  IV  NOT_4285(g21070,I20937);
  IV  NOT_4286(g6888,I11701);
  IV  NOT_4287(g22974,g20330);
  IV  NOT_4288(g32831,g31376);
  IV  NOT_4289(g33691,I31528);
  IV  NOT_4290(g32445,I29973);
  IV  NOT_4291(I32938,g34663);
  IV  NOT_4292(I32093,g33670);
  IV  NOT_4293(I13276,g5798);
  IV  NOT_4294(g16716,g13948);
  IV  NOT_4295(g9678,g5406);
  IV  NOT_4296(g10039,g2273);
  IV  NOT_4297(g10306,I13726);
  IV  NOT_4298(g32499,g31376);
  IV  NOT_4299(g23986,g18833);
  IV  NOT_4300(g30591,I28851);
  IV  NOT_4301(g6956,g4242);
  IV  NOT_4302(g18984,g17486);
  IV  NOT_4303(g8623,g3990);
  IV  NOT_4304(I11809,g6741);
  IV  NOT_4305(g34591,I32681);
  IV  NOT_4306(I18214,g12918);
  IV  NOT_4307(g12892,g10398);
  IV  NOT_4308(g34785,I32985);
  IV  NOT_4309(g16582,g13915);
  IV  NOT_4310(g17772,g14297);
  IV  NOT_4311(g34776,I32970);
  IV  NOT_4312(g11425,g7640);
  IV  NOT_4313(g10038,g2241);
  IV  NOT_4314(g32498,g31566);
  IV  NOT_4315(g23384,I22485);
  IV  NOT_4316(g17639,I18600);
  IV  NOT_4317(I12141,g599);
  IV  NOT_4318(g34147,g33823);
  IV  NOT_4319(g9682,I13280);
  IV  NOT_4320(g9766,g2748);
  IV  NOT_4321(g15811,g13125);
  IV  NOT_4322(g16310,g13223);
  IV  NOT_4323(g7096,g6537);
  IV  NOT_4324(g10815,g9917);
  IV  NOT_4325(g13458,g11048);
  IV  NOT_4326(g24160,I23324);
  IV  NOT_4327(I15918,g12381);
  IV  NOT_4328(g9305,g5381);
  IV  NOT_4329(g7496,g5969);
  IV  NOT_4330(g33929,I31803);
  IV  NOT_4331(g16627,I17819);
  IV  NOT_4332(g17638,g14838);
  IV  NOT_4333(g22841,g20391);
  IV  NOT_4334(g34950,g34940);
  IV  NOT_4335(g12914,g12235);
  IV  NOT_4336(g13010,I15620);
  IV  NOT_4337(g32611,g31154);
  IV  NOT_4338(g7845,g1146);
  IV  NOT_4339(I33232,g34957);
  IV  NOT_4340(g25451,g22228);
  IV  NOT_4341(g32722,g30937);
  IV  NOT_4342(g25220,I24396);
  IV  NOT_4343(g32924,g30937);
  IV  NOT_4344(g33928,I31800);
  IV  NOT_4345(g19947,g17226);
  IV  NOT_4346(g7195,g25);
  IV  NOT_4347(g12907,g10415);
  IV  NOT_4348(g20617,g15277);
  IV  NOT_4349(g17416,g14956);
  IV  NOT_4350(g7395,g6005);
  IV  NOT_4351(g7891,g2994);
  IV  NOT_4352(g8651,g758);
  IV  NOT_4353(g16958,g14238);
  IV  NOT_4354(g9748,g114);
  IV  NOT_4355(g13545,I16010);
  IV  NOT_4356(g23877,g19147);
  IV  NOT_4357(g19273,g16100);
  IV  NOT_4358(g20915,I20882);
  IV  NOT_4359(g7913,g1052);
  IV  NOT_4360(g27074,I25790);
  IV  NOT_4361(g28321,g27317);
  IV  NOT_4362(I32837,g34498);
  IV  NOT_4363(g30996,g29694);
  IV  NOT_4364(g25246,g23828);
  IV  NOT_4365(g34151,I32106);
  IV  NOT_4366(I12135,g807);
  IV  NOT_4367(g10143,g568);
  IV  NOT_4368(g29213,I27555);
  IV  NOT_4369(g34996,I33288);
  IV  NOT_4370(g23019,g19866);
  IV  NOT_4371(I33261,g34977);
  IV  NOT_4372(g8285,I12497);
  IV  NOT_4373(g12074,I14932);
  IV  NOT_4374(I25695,g25690);
  IV  NOT_4375(g9226,g1564);
  IV  NOT_4376(g20277,g16487);
  IV  NOT_4377(g16603,I17787);
  IV  NOT_4378(g16742,g13983);
  IV  NOT_4379(g23196,g20785);
  IV  NOT_4380(g34844,g34737);
  IV  NOT_4381(I22564,g20857);
  IV  NOT_4382(g16096,g13530);
  IV  NOT_4383(g23018,g19801);
  IV  NOT_4384(g32753,g30735);
  IV  NOT_4385(g12238,I15102);
  IV  NOT_4386(g32461,g30614);
  IV  NOT_4387(I21242,g16540);
  IV  NOT_4388(g10169,g6395);
  IV  NOT_4389(g24075,g19935);
  IV  NOT_4390(g17579,g14959);
  IV  NOT_4391(g19371,I19857);
  IV  NOT_4392(g20595,g15877);
  IV  NOT_4393(g23526,g21611);
  IV  NOT_4394(g6808,g554);
  IV  NOT_4395(g20494,g17847);
  IV  NOT_4396(g14169,g12381);
  IV  NOT_4397(g8139,g1648);
  IV  NOT_4398(I16289,g12107);
  IV  NOT_4399(I32455,g34242);
  IV  NOT_4400(g7266,g35);
  IV  NOT_4401(g29912,g28827);
  IV  NOT_4402(g29311,g28998);
  IV  NOT_4403(g10410,g7069);
  IV  NOT_4404(g20623,g17929);
  IV  NOT_4405(g27675,I26309);
  IV  NOT_4406(I12049,g781);
  IV  NOT_4407(g9373,g5142);
  IV  NOT_4408(g17014,g14297);
  IV  NOT_4409(g27092,g26737);
  IV  NOT_4410(g9091,g1430);
  IV  NOT_4411(g20037,g17328);
  IV  NOT_4412(g31827,g29385);
  IV  NOT_4413(g32736,g30937);
  IV  NOT_4414(I32617,g34333);
  IV  NOT_4415(g13322,g10918);
  IV  NOT_4416(g32887,g30614);
  IV  NOT_4417(I32470,g34247);
  IV  NOT_4418(g24623,g23076);
  IV  NOT_4419(g33827,I31672);
  IV  NOT_4420(g9491,g2729);
  IV  NOT_4421(I14905,g9822);
  IV  NOT_4422(g24037,g21127);
  IV  NOT_4423(g34420,g34152);
  IV  NOT_4424(g16429,I17671);
  IV  NOT_4425(I11665,g1589);
  IV  NOT_4426(g20782,g15853);
  IV  NOT_4427(g21457,g17367);
  IV  NOT_4428(g13901,g11480);
  IV  NOT_4429(g23402,g20875);
  IV  NOT_4430(I13166,g5101);
  IV  NOT_4431(g32529,g30735);
  IV  NOT_4432(g23457,I22580);
  IV  NOT_4433(g25370,g22228);
  IV  NOT_4434(g8795,I12793);
  IV  NOT_4435(g10363,I13779);
  IV  NOT_4436(I24400,g23954);
  IV  NOT_4437(g10217,g2102);
  IV  NOT_4438(I14593,g9978);
  IV  NOT_4439(g30318,g28274);
  IV  NOT_4440(g14363,I16521);
  IV  NOT_4441(g14217,I16417);
  IV  NOT_4442(g9283,g1736);
  IV  NOT_4443(I14346,g10233);
  IV  NOT_4444(g16428,I17668);
  IV  NOT_4445(g9369,g5084);
  IV  NOT_4446(g32528,g31554);
  IV  NOT_4447(g32696,g30825);
  IV  NOT_4448(g9007,g1083);
  IV  NOT_4449(I21230,g16540);
  IV  NOT_4450(g32843,g31021);
  IV  NOT_4451(g6957,g2932);
  IV  NOT_4452(g24419,g22722);
  IV  NOT_4453(g32393,g30922);
  IV  NOT_4454(g9407,g6549);
  IV  NOT_4455(I15295,g8515);
  IV  NOT_4456(I11892,g4408);
  IV  NOT_4457(g34059,g33658);
  IV  NOT_4458(g8672,g4669);
  IV  NOT_4459(g9920,g4322);
  IV  NOT_4460(I15144,g5659);
  IV  NOT_4461(I13892,g1576);
  IV  NOT_4462(g31803,g29385);
  IV  NOT_4463(g32764,g30937);
  IV  NOT_4464(g24155,I23309);
  IV  NOT_4465(g24418,g22722);
  IV  NOT_4466(I32467,g34246);
  IV  NOT_4467(g20266,g17873);
  IV  NOT_4468(g8477,g3061);
  IV  NOT_4469(g34540,I32607);
  IV  NOT_4470(g11823,I14647);
  IV  NOT_4471(g13680,I16077);
  IV  NOT_4472(g17615,I18574);
  IV  NOT_4473(g12883,g10390);
  IV  NOT_4474(g13144,I15773);
  IV  NOT_4475(g22493,g19801);
  IV  NOT_4476(g7097,I11809);
  IV  NOT_4477(g23001,g19801);
  IV  NOT_4478(g34058,g33660);
  IV  NOT_4479(g24170,I23354);
  IV  NOT_4480(g32869,g30735);
  IV  NOT_4481(I18882,g16580);
  IV  NOT_4482(g32960,g31327);
  IV  NOT_4483(I18414,g14359);
  IV  NOT_4484(g7497,g6358);
  IV  NOT_4485(I14797,g9636);
  IV  NOT_4486(g19421,g16326);
  IV  NOT_4487(g17720,g15045);
  IV  NOT_4488(I33056,g34778);
  IV  NOT_4489(I25689,g25688);
  IV  NOT_4490(g9582,g703);
  IV  NOT_4491(g11336,g7620);
  IV  NOT_4492(g7960,g1404);
  IV  NOT_4493(g32868,g31376);
  IV  NOT_4494(g8205,g2208);
  IV  NOT_4495(I32782,g34571);
  IV  NOT_4496(g10223,g4561);
  IV  NOT_4497(g21689,I21250);
  IV  NOT_4498(g23256,g20785);
  IV  NOT_4499(I12106,g626);
  IV  NOT_4500(I12605,g1570);
  IV  NOT_4501(g17430,I18373);
  IV  NOT_4502(g17746,g14825);
  IV  NOT_4503(g20853,g15595);
  IV  NOT_4504(g34044,g33675);
  IV  NOT_4505(g21280,g16601);
  IV  NOT_4506(g23923,g18997);
  IV  NOT_4507(I14409,g8364);
  IV  NOT_4508(g29152,g27907);
  IV  NOT_4509(g29846,g28391);
  IV  NOT_4510(I32352,g34169);
  IV  NOT_4511(I29002,g29675);
  IV  NOT_4512(g21300,I21047);
  IV  NOT_4513(g20167,g16971);
  IV  NOT_4514(g20194,g16897);
  IV  NOT_4515(g20589,g15224);
  IV  NOT_4516(g32709,g30735);
  IV  NOT_4517(g11966,I14800);
  IV  NOT_4518(g23300,g20283);
  IV  NOT_4519(I12463,g4812);
  IV  NOT_4520(g17465,g12955);
  IV  NOT_4521(g8742,g4035);
  IV  NOT_4522(g13966,I16246);
  IV  NOT_4523(g10084,g2837);
  IV  NOT_4524(g24167,I23345);
  IV  NOT_4525(g9415,g2169);
  IV  NOT_4526(g19541,g16136);
  IV  NOT_4527(g30301,I28548);
  IV  NOT_4528(g10110,g661);
  IV  NOT_4529(g11631,g8595);
  IV  NOT_4530(g19473,g16349);
  IV  NOT_4531(g18101,I18909);
  IV  NOT_4532(g11017,g10289);
  IV  NOT_4533(g20588,g18008);
  IV  NOT_4534(g20524,g17873);
  IV  NOT_4535(g32708,g31376);
  IV  NOT_4536(I32170,g33638);
  IV  NOT_4537(I12033,g776);
  IV  NOT_4538(g13017,I15633);
  IV  NOT_4539(I28174,g28803);
  IV  NOT_4540(I29245,g29491);
  IV  NOT_4541(g32471,g31376);
  IV  NOT_4542(g19789,g17015);
  IV  NOT_4543(g24524,g22876);
  IV  NOT_4544(g24836,I24008);
  IV  NOT_4545(g16129,I17488);
  IV  NOT_4546(g25227,g22763);
  IV  NOT_4547(g14321,g10874);
  IV  NOT_4548(g34739,I32909);
  IV  NOT_4549(g10531,g8925);
  IV  NOT_4550(g17684,g15036);
  IV  NOT_4551(g27438,I26130);
  IV  NOT_4552(g14179,g11048);
  IV  NOT_4553(g25025,g22498);
  IV  NOT_4554(g7267,g1604);
  IV  NOT_4555(g24477,I23680);
  IV  NOT_4556(g10178,g2126);
  IV  NOT_4557(g26632,g25473);
  IV  NOT_4558(g24119,g19935);
  IV  NOT_4559(g27349,g26352);
  IV  NOT_4560(I31650,g33212);
  IV  NOT_4561(g23066,g20330);
  IV  NOT_4562(I28390,g29185);
  IV  NOT_4563(g9721,g5097);
  IV  NOT_4564(g23231,g20050);
  IV  NOT_4565(g34699,I32855);
  IV  NOT_4566(g19434,g16326);
  IV  NOT_4567(g16626,g14133);
  IV  NOT_4568(g8273,g2453);
  IV  NOT_4569(g10685,I13995);
  IV  NOT_4570(I16489,g12793);
  IV  NOT_4571(g16323,I17653);
  IV  NOT_4572(g24118,g19890);
  IV  NOT_4573(g10373,g6917);
  IV  NOT_4574(g14186,g11346);
  IV  NOT_4575(g14676,I16775);
  IV  NOT_4576(g24022,g20982);
  IV  NOT_4577(g34698,g34550);
  IV  NOT_4578(g7293,g4452);
  IV  NOT_4579(g12906,g10413);
  IV  NOT_4580(g16533,I17733);
  IV  NOT_4581(g20616,g15277);
  IV  NOT_4582(I18114,g14509);
  IV  NOT_4583(g23876,g19074);
  IV  NOT_4584(I18758,g6719);
  IV  NOT_4585(g13023,g11897);
  IV  NOT_4586(g18874,g15938);
  IV  NOT_4587(I31528,g33219);
  IV  NOT_4588(g25044,g23675);
  IV  NOT_4589(I19661,g17587);
  IV  NOT_4590(g29929,g28914);
  IV  NOT_4591(g16775,I17999);
  IV  NOT_4592(I18107,g4019);
  IV  NOT_4593(g10417,g7117);
  IV  NOT_4594(I25511,g25073);
  IV  NOT_4595(g32602,g30825);
  IV  NOT_4596(g32810,g31376);
  IV  NOT_4597(I13637,g102);
  IV  NOT_4598(I20882,g17619);
  IV  NOT_4599(g32657,g31528);
  IV  NOT_4600(g32774,g30735);
  IV  NOT_4601(g33778,I31625);
  IV  NOT_4602(g7828,g4871);
  IV  NOT_4603(g32955,g30735);
  IV  NOT_4604(g21511,g15483);
  IV  NOT_4605(g29928,g28871);
  IV  NOT_4606(I26670,g27709);
  IV  NOT_4607(g20704,g15373);
  IV  NOT_4608(g23511,I22640);
  IV  NOT_4609(g34427,I32452);
  IV  NOT_4610(I32119,g33648);
  IV  NOT_4611(g32879,g31327);
  IV  NOT_4612(g8572,I12654);
  IV  NOT_4613(g20053,g17328);
  IV  NOT_4614(g32970,g30825);
  IV  NOT_4615(g10334,g4420);
  IV  NOT_4616(g19682,g17015);
  IV  NOT_4617(I14537,g10106);
  IV  NOT_4618(g24053,g21256);
  IV  NOT_4619(g25120,g22432);
  IV  NOT_4620(I17780,g13303);
  IV  NOT_4621(g17523,g14732);
  IV  NOT_4622(g20900,I20864);
  IV  NOT_4623(g8712,I12712);
  IV  NOT_4624(g7592,g347);
  IV  NOT_4625(I16544,g11931);
  IV  NOT_4626(I18849,g14290);
  IV  NOT_4627(g18008,I18868);
  IV  NOT_4628(g32878,g30937);
  IV  NOT_4629(g31945,g31189);
  IV  NOT_4630(g21660,g17694);
  IV  NOT_4631(g24466,I23671);
  IV  NOT_4632(I16713,g5331);
  IV  NOT_4633(g9689,g124);
  IV  NOT_4634(g10762,g8470);
  IV  NOT_4635(g25562,g22763);
  IV  NOT_4636(g18892,g15680);
  IV  NOT_4637(g20036,g17433);
  IV  NOT_4638(g31826,g29385);
  IV  NOT_4639(g32886,g31327);
  IV  NOT_4640(I33161,g34894);
  IV  NOT_4641(I18398,g13745);
  IV  NOT_4642(g20101,g17533);
  IV  NOT_4643(g24036,g20982);
  IV  NOT_4644(I12541,g194);
  IV  NOT_4645(g20560,g17328);
  IV  NOT_4646(g16856,I18048);
  IV  NOT_4647(g21456,g15509);
  IV  NOT_4648(I26667,g27585);
  IV  NOT_4649(g11985,I14827);
  IV  NOT_4650(g17475,I18398);
  IV  NOT_4651(g24101,g20998);
  IV  NOT_4652(I23684,g23230);
  IV  NOT_4653(g32792,g31710);
  IV  NOT_4654(g23456,g21514);
  IV  NOT_4655(g13976,g11130);
  IV  NOT_4656(g24177,I23375);
  IV  NOT_4657(g24560,g22942);
  IV  NOT_4658(I15954,g12381);
  IV  NOT_4659(g32967,g31327);
  IV  NOT_4660(g10216,I13684);
  IV  NOT_4661(g14423,I16579);
  IV  NOT_4662(g8534,g3338);
  IV  NOT_4663(I16610,g10981);
  IV  NOT_4664(g9671,g5134);
  IV  NOT_4665(g20642,g15277);
  IV  NOT_4666(g23480,I22601);
  IV  NOT_4667(g27415,g26382);
  IV  NOT_4668(I20584,g16587);
  IV  NOT_4669(g23916,g19277);
  IV  NOT_4670(g9030,g4793);
  IV  NOT_4671(g19760,g17015);
  IV  NOT_4672(I32305,g34209);
  IV  NOT_4673(I14381,g8300);
  IV  NOT_4674(g16512,g14015);
  IV  NOT_4675(I16679,g12039);
  IV  NOT_4676(g23550,g20248);
  IV  NOT_4677(g26784,g25341);
  IV  NOT_4678(g9247,g1559);
  IV  NOT_4679(I33258,g34976);
  IV  NOT_4680(I32809,g34586);
  IV  NOT_4681(g18907,g15979);
  IV  NOT_4682(g7624,I12106);
  IV  NOT_4683(g32459,g31070);
  IV  NOT_4684(g20064,g17533);
  IV  NOT_4685(g7953,g4966);
  IV  NOT_4686(g30572,g29945);
  IV  NOT_4687(g24064,g20841);
  IV  NOT_4688(g28579,g27714);
  IV  NOT_4689(g9564,g6120);
  IV  NOT_4690(I18135,g13144);
  IV  NOT_4691(g23307,g20924);
  IV  NOT_4692(g32919,g30735);
  IV  NOT_4693(g23085,g19957);
  IV  NOT_4694(g32458,g30825);
  IV  NOT_4695(I24759,g24229);
  IV  NOT_4696(g14543,I16660);
  IV  NOT_4697(g33932,I31810);
  IV  NOT_4698(g9826,g1844);
  IV  NOT_4699(g10117,g2509);
  IV  NOT_4700(g10000,g6151);
  IV  NOT_4701(g26824,g25298);
  IV  NOT_4702(I16460,g10430);
  IV  NOT_4703(g20874,g15680);
  IV  NOT_4704(g21054,g15373);
  IV  NOT_4705(g32918,g31327);
  IV  NOT_4706(g23243,g21070);
  IV  NOT_4707(g20630,g17955);
  IV  NOT_4708(g11842,I14660);
  IV  NOT_4709(g21431,g18065);
  IV  NOT_4710(g9741,I13317);
  IV  NOT_4711(g8903,g1075);
  IV  NOT_4712(g23431,g21514);
  IV  NOT_4713(I13906,g7620);
  IV  NOT_4714(g32545,g31070);
  IV  NOT_4715(g9910,g2108);
  IV  NOT_4716(g17600,g14659);
  IV  NOT_4717(I19671,g15932);
  IV  NOT_4718(g34490,I32547);
  IV  NOT_4719(g20166,g16886);
  IV  NOT_4720(g20009,g16349);
  IV  NOT_4721(I22583,g20998);
  IV  NOT_4722(g27576,g26081);
  IV  NOT_4723(g27585,g25994);
  IV  NOT_4724(g20665,g15373);
  IV  NOT_4725(g25547,g22550);
  IV  NOT_4726(g32599,g30673);
  IV  NOT_4727(I20744,g17141);
  IV  NOT_4728(I31810,g33164);
  IV  NOT_4729(g9638,g1620);
  IV  NOT_4730(g21269,g15506);
  IV  NOT_4731(g24166,I23342);
  IV  NOT_4732(g24665,g23067);
  IV  NOT_4733(g7716,g1199);
  IV  NOT_4734(g7149,g4564);
  IV  NOT_4735(g34784,I32982);
  IV  NOT_4736(g7349,g1270);
  IV  NOT_4737(g30297,g28758);
  IV  NOT_4738(g27554,g26625);
  IV  NOT_4739(g20008,g16449);
  IV  NOT_4740(g34956,I33214);
  IV  NOT_4741(g17952,I18858);
  IV  NOT_4742(g32598,g30614);
  IV  NOT_4743(g13016,g11878);
  IV  NOT_4744(I22046,g19330);
  IV  NOT_4745(g23942,g21562);
  IV  NOT_4746(I20399,g16205);
  IV  NOT_4747(g23341,g21163);
  IV  NOT_4748(g18092,I18882);
  IV  NOT_4749(g21268,g15680);
  IV  NOT_4750(I14192,g10233);
  IV  NOT_4751(I18048,g13638);
  IV  NOT_4752(I28062,g29194);
  IV  NOT_4753(g25226,g22763);
  IV  NOT_4754(g22137,g21370);
  IV  NOT_4755(g21156,g17247);
  IV  NOT_4756(g17821,I18829);
  IV  NOT_4757(g8178,I12437);
  IV  NOT_4758(g6801,g391);
  IV  NOT_4759(I21006,g15579);
  IV  NOT_4760(g28615,g27817);
  IV  NOT_4761(I16875,g6675);
  IV  NOT_4762(g25481,g22228);
  IV  NOT_4763(I15893,g10430);
  IV  NOT_4764(I31878,g33696);
  IV  NOT_4765(g19649,g17015);
  IV  NOT_4766(I32874,g34504);
  IV  NOT_4767(g21180,g18008);
  IV  NOT_4768(I14663,g9747);
  IV  NOT_4769(g21670,g16540);
  IV  NOT_4770(I18221,g13605);
  IV  NOT_4771(g16722,I17938);
  IV  NOT_4772(g16924,I18092);
  IV  NOT_4773(g20555,g15480);
  IV  NOT_4774(g32817,g31376);
  IV  NOT_4775(I28851,g29317);
  IV  NOT_4776(I28872,g30072);
  IV  NOT_4777(I32693,g34433);
  IV  NOT_4778(g8135,I12418);
  IV  NOT_4779(I21222,g18091);
  IV  NOT_4780(g19491,g16349);
  IV  NOT_4781(g34181,g33913);
  IV  NOT_4782(g34671,I32797);
  IV  NOT_4783(g20570,g15277);
  IV  NOT_4784(g20712,g15509);
  IV  NOT_4785(g11865,g10124);
  IV  NOT_4786(I22302,g19353);
  IV  NOT_4787(g13865,I16168);
  IV  NOT_4788(g20914,g15373);
  IV  NOT_4789(g21335,I21067);
  IV  NOT_4790(g18883,g15938);
  IV  NOT_4791(g32532,g31170);
  IV  NOT_4792(g32901,g31327);
  IV  NOT_4793(g14639,I16747);
  IV  NOT_4794(g10230,I13694);
  IV  NOT_4795(g23335,g20391);
  IV  NOT_4796(I32665,g34386);
  IV  NOT_4797(g19755,g15915);
  IV  NOT_4798(g6755,I11620);
  IV  NOT_4799(g12921,g12228);
  IV  NOT_4800(g23839,g18997);
  IV  NOT_4801(I17787,g3267);
  IV  NOT_4802(g17873,I18849);
  IV  NOT_4803(g23930,g19147);
  IV  NOT_4804(g23993,g19277);
  IV  NOT_4805(g32783,g30825);
  IV  NOT_4806(g19770,g17062);
  IV  NOT_4807(I29199,g30237);
  IV  NOT_4808(g30931,I28913);
  IV  NOT_4809(g8805,I12799);
  IV  NOT_4810(I14862,g8092);
  IV  NOT_4811(g8916,I12887);
  IV  NOT_4812(I16160,g11237);
  IV  NOT_4813(g21694,g16540);
  IV  NOT_4814(g23838,g18997);
  IV  NOT_4815(g9861,g5459);
  IV  NOT_4816(g10416,g10318);
  IV  NOT_4817(I15705,g12218);
  IV  NOT_4818(g9048,I12963);
  IV  NOT_4819(I17302,g14044);
  IV  NOT_4820(g32561,g30614);
  IV  NOT_4821(g32656,g30673);
  IV  NOT_4822(g23965,g21611);
  IV  NOT_4823(I31459,g33219);
  IV  NOT_4824(g20239,g17128);
  IV  NOT_4825(I32476,g34277);
  IV  NOT_4826(g11705,I14576);
  IV  NOT_4827(I22640,g21256);
  IV  NOT_4828(g24074,g21193);
  IV  NOT_4829(I22769,g21277);
  IV  NOT_4830(g26860,I25594);
  IV  NOT_4831(I14326,g8607);
  IV  NOT_4832(g34426,I32449);
  IV  NOT_4833(g11042,g8691);
  IV  NOT_4834(g16031,I17436);
  IV  NOT_4835(g20567,g15426);
  IV  NOT_4836(g20594,g15277);
  IV  NOT_4837(g32680,g31376);
  IV  NOT_4838(g10391,g6988);
  IV  NOT_4839(I16455,g11845);
  IV  NOT_4840(g32823,g31327);
  IV  NOT_4841(g20238,g17096);
  IV  NOT_4842(g25297,g23746);
  IV  NOT_4843(g13255,g10632);
  IV  NOT_4844(g9827,g1974);
  IV  NOT_4845(g13189,g10762);
  IV  NOT_4846(g22542,g19801);
  IV  NOT_4847(g13679,g10573);
  IV  NOT_4848(g28142,I26649);
  IV  NOT_4849(g31811,g29385);
  IV  NOT_4850(g23487,g20924);
  IV  NOT_4851(g14510,I16629);
  IV  NOT_4852(g31646,I29228);
  IV  NOT_4853(g9333,g417);
  IV  NOT_4854(I14702,g7717);
  IV  NOT_4855(g19794,g16489);
  IV  NOT_4856(g11678,I14563);
  IV  NOT_4857(g12184,I15036);
  IV  NOT_4858(g16529,g14055);
  IV  NOT_4859(g29081,g27837);
  IV  NOT_4860(g12805,g9511);
  IV  NOT_4861(g13188,g10909);
  IV  NOT_4862(g19395,g16431);
  IV  NOT_4863(g23502,g21070);
  IV  NOT_4864(I27927,g28803);
  IV  NOT_4865(g20382,g15171);
  IV  NOT_4866(I16201,g4023);
  IV  NOT_4867(I23351,g23263);
  IV  NOT_4868(I31545,g33219);
  IV  NOT_4869(I23372,g23361);
  IV  NOT_4870(g26700,g25429);
  IV  NOT_4871(g7258,g4414);
  IV  NOT_4872(I33079,g34809);
  IV  NOT_4873(g11686,I14567);
  IV  NOT_4874(g16528,g14154);
  IV  NOT_4875(g7577,g1263);
  IV  NOT_4876(g7867,g1489);
  IV  NOT_4877(g13460,I15942);
  IV  NOT_4878(g15831,g13385);
  IV  NOT_4879(I26479,g25771);
  IV  NOT_4880(I12927,g4332);
  IV  NOT_4881(g26987,g26131);
  IV  NOT_4882(g11383,g9061);
  IV  NOT_4883(g10014,g6439);
  IV  NOT_4884(g23443,g21468);
  IV  NOT_4885(I15030,g10073);
  IV  NOT_4886(I18795,g5327);
  IV  NOT_4887(g21279,g15680);
  IV  NOT_4888(g24176,I23372);
  IV  NOT_4889(g24185,I23399);
  IV  NOT_4890(g23279,g21037);
  IV  NOT_4891(g32966,g31021);
  IV  NOT_4892(g19633,g16931);
  IV  NOT_4893(g7717,I12172);
  IV  NOT_4894(g30088,g29094);
  IV  NOT_4895(g24092,g20857);
  IV  NOT_4896(I32074,g33670);
  IV  NOT_4897(g29945,I28174);
  IV  NOT_4898(g6868,I11688);
  IV  NOT_4899(g11030,g8292);
  IV  NOT_4900(g20154,I20412);
  IV  NOT_4901(g22905,I22114);
  IV  NOT_4902(g32631,g30825);
  IV  NOT_4903(g19719,g16897);
  IV  NOT_4904(g21278,I21013);
  IV  NOT_4905(g11294,g7598);
  IV  NOT_4906(g24154,I23306);
  IV  NOT_4907(I32594,g34298);
  IV  NOT_4908(g8037,g405);
  IV  NOT_4909(g23278,g20283);
  IV  NOT_4910(g13267,I15831);
  IV  NOT_4911(g29999,g28973);
  IV  NOT_4912(g32364,I29894);
  IV  NOT_4913(g6767,I11626);
  IV  NOT_4914(g17614,I18571);
  IV  NOT_4915(g22593,g19801);
  IV  NOT_4916(g9780,I13360);
  IV  NOT_4917(g16960,I18114);
  IV  NOT_4918(g20637,g15224);
  IV  NOT_4919(g26943,I25695);
  IV  NOT_4920(g8102,g3072);
  IV  NOT_4921(g13065,g10476);
  IV  NOT_4922(g19718,g17015);
  IV  NOT_4923(g21286,g15509);
  IV  NOT_4924(g8302,g1926);
  IV  NOT_4925(g14442,I16593);
  IV  NOT_4926(g29998,g28966);
  IV  NOT_4927(g17607,I18560);
  IV  NOT_4928(g21468,I21181);
  IV  NOT_4929(g17320,I18297);
  IV  NOT_4930(g21306,g15582);
  IV  NOT_4931(g31850,g29385);
  IV  NOT_4932(g8579,g2771);
  IV  NOT_4933(g23306,g20924);
  IV  NOT_4934(I29225,g30311);
  IV  NOT_4935(I31817,g33323);
  IV  NOT_4936(g7975,g3040);
  IV  NOT_4937(g33850,I31701);
  IV  NOT_4938(g17530,g14947);
  IV  NOT_4939(g10116,g2413);
  IV  NOT_4940(g9662,g3983);
  IV  NOT_4941(g9018,g4273);
  IV  NOT_4942(g11875,I14687);
  IV  NOT_4943(g8719,I12719);
  IV  NOT_4944(g27013,I25743);
  IV  NOT_4945(g7026,g5507);
  IV  NOT_4946(I32675,g34427);
  IV  NOT_4947(g9467,g6434);
  IV  NOT_4948(g19440,g15915);
  IV  NOT_4949(g16709,I17919);
  IV  NOT_4950(g17122,g14348);
  IV  NOT_4951(g34126,I32067);
  IV  NOT_4952(g34659,I32775);
  IV  NOT_4953(I12770,g4200);
  IV  NOT_4954(I12563,g3798);
  IV  NOT_4955(g12013,I14866);
  IV  NOT_4956(g23815,g19074);
  IV  NOT_4957(g34987,I33261);
  IV  NOT_4958(I25677,g25640);
  IV  NOT_4959(I15837,g1459);
  IV  NOT_4960(I33158,g34897);
  IV  NOT_4961(g7170,g5719);
  IV  NOT_4962(g19861,g17096);
  IV  NOT_4963(g10275,g4584);
  IV  NOT_4964(g19573,g16877);
  IV  NOT_4965(g8917,I12890);
  IV  NOT_4966(g16708,I17916);
  IV  NOT_4967(g22153,g18997);
  IV  NOT_4968(g21677,I21238);
  IV  NOT_4969(g33228,I30766);
  IV  NOT_4970(g10430,I13847);
  IV  NOT_4971(g14275,g12358);
  IV  NOT_4972(g25546,g22550);
  IV  NOT_4973(g32571,g31376);
  IV  NOT_4974(I31561,g33197);
  IV  NOT_4975(I17249,g13605);
  IV  NOT_4976(g25211,g22763);
  IV  NOT_4977(I32935,g34657);
  IV  NOT_4978(g22409,I21860);
  IV  NOT_4979(g19389,g17532);
  IV  NOT_4980(g17641,g14845);
  IV  NOT_4981(g20501,g17955);
  IV  NOT_4982(g26870,I25606);
  IV  NOT_4983(g30296,g28889);
  IV  NOT_4984(g20577,g15483);
  IV  NOT_4985(g34339,g34077);
  IV  NOT_4986(g9816,g6167);
  IV  NOT_4987(g34943,I33197);
  IV  NOT_4988(I20951,g17782);
  IV  NOT_4989(g25024,g22472);
  IV  NOT_4990(g33716,I31569);
  IV  NOT_4991(I31823,g33149);
  IV  NOT_4992(g19612,g16897);
  IV  NOT_4993(g34296,I32297);
  IV  NOT_4994(g7280,g2153);
  IV  NOT_4995(g29897,I28128);
  IV  NOT_4996(g7939,g1280);
  IV  NOT_4997(g22136,g20277);
  IV  NOT_4998(g29961,g28892);
  IV  NOT_4999(g8442,g3476);
  IV  NOT_5000(g22408,g19483);
  IV  NOT_5001(g22635,g19801);
  IV  NOT_5002(I12767,g4197);
  IV  NOT_5003(g14237,g11666);
  IV  NOT_5004(g8786,I12770);
  IV  NOT_5005(g23937,g19277);
  IV  NOT_5006(g10035,g1720);
  IV  NOT_5007(g32495,g31070);
  IV  NOT_5008(g29505,g29186);
  IV  NOT_5009(g19777,g17015);
  IV  NOT_5010(g17409,I18344);
  IV  NOT_5011(I12899,g4232);
  IV  NOT_5012(g7544,g918);
  IV  NOT_5013(g8164,g3484);
  IV  NOT_5014(g9381,g5527);
  IV  NOT_5015(I15617,g12037);
  IV  NOT_5016(I13805,g6976);
  IV  NOT_5017(I18788,g13138);
  IV  NOT_5018(g8364,g1585);
  IV  NOT_5019(g32816,g31327);
  IV  NOT_5020(I15915,g10430);
  IV  NOT_5021(g24438,g22722);
  IV  NOT_5022(g11470,g7625);
  IV  NOT_5023(g17136,g14348);
  IV  NOT_5024(g10142,I13637);
  IV  NOT_5025(g17408,I18341);
  IV  NOT_5026(g34060,g33704);
  IV  NOT_5027(g29212,I27552);
  IV  NOT_5028(g7636,g4098);
  IV  NOT_5029(g9685,g6533);
  IV  NOT_5030(I26676,g27736);
  IV  NOT_5031(g9197,g1221);
  IV  NOT_5032(I18829,g13350);
  IV  NOT_5033(g32687,g31376);
  IV  NOT_5034(g9397,g6088);
  IV  NOT_5035(I18434,g13782);
  IV  NOT_5036(g33959,I31878);
  IV  NOT_5037(g9021,I12954);
  IV  NOT_5038(I12719,g365);
  IV  NOT_5039(g16602,g14101);
  IV  NOT_5040(g21410,g15224);
  IV  NOT_5041(g34197,g33812);
  IV  NOT_5042(I27718,g28231);
  IV  NOT_5043(I16401,g869);
  IV  NOT_5044(g16774,g14024);
  IV  NOT_5045(g23410,g21562);
  IV  NOT_5046(g8770,g749);
  IV  NOT_5047(I29337,g30286);
  IV  NOT_5048(g34855,I33079);
  IV  NOT_5049(I26654,g27576);
  IV  NOT_5050(I22380,g21156);
  IV  NOT_5051(g16955,I18107);
  IV  NOT_5052(g32752,g31376);
  IV  NOT_5053(g8296,g246);
  IV  NOT_5054(g25250,I24434);
  IV  NOT_5055(g27100,g26759);
  IV  NOT_5056(g32954,g31376);
  IV  NOT_5057(g8725,g739);
  IV  NOT_5058(g24083,g19984);
  IV  NOT_5059(g33378,I30904);
  IV  NOT_5060(g21666,g16540);
  IV  NOT_5061(g23479,g21562);
  IV  NOT_5062(I26936,g27599);
  IV  NOT_5063(g32643,g31376);
  IV  NOT_5064(g6940,g4035);
  IV  NOT_5065(I15494,g10385);
  IV  NOT_5066(g13075,I15705);
  IV  NOT_5067(g23363,I22470);
  IV  NOT_5068(I18344,g13003);
  IV  NOT_5069(g7187,g6065);
  IV  NOT_5070(g7387,g2421);
  IV  NOT_5071(g20622,g15595);
  IV  NOT_5072(g11467,g7623);
  IV  NOT_5073(g13595,g10951);
  IV  NOT_5074(I17999,g4012);
  IV  NOT_5075(g20566,g15224);
  IV  NOT_5076(g7461,g2567);
  IV  NOT_5077(I15623,g12040);
  IV  NOT_5078(g23478,g21514);
  IV  NOT_5079(g13494,g11912);
  IV  NOT_5080(g23015,g20391);
  IV  NOT_5081(g8553,g3747);
  IV  NOT_5082(I26334,g26834);
  IV  NOT_5083(I19707,g17590);
  IV  NOT_5084(g25296,g23745);
  IV  NOT_5085(g10130,g5694);
  IV  NOT_5086(g16171,g13530);
  IV  NOT_5087(g33944,I31829);
  IV  NOT_5088(g19061,I19762);
  IV  NOT_5089(g26818,I25530);
  IV  NOT_5090(g16886,I18078);
  IV  NOT_5091(I27573,g28157);
  IV  NOT_5092(g32669,g30614);
  IV  NOT_5093(I15782,g10430);
  IV  NOT_5094(g23486,g20785);
  IV  NOT_5095(g26055,I25115);
  IV  NOT_5096(g13037,g10981);
  IV  NOT_5097(g10362,g6850);
  IV  NOT_5098(g29149,g27837);
  IV  NOT_5099(g7027,g5499);
  IV  NOT_5100(I19818,g1056);
  IV  NOT_5101(g19766,g16449);
  IV  NOT_5102(g21556,g15669);
  IV  NOT_5103(I12861,g4372);
  IV  NOT_5104(g10165,g5698);
  IV  NOT_5105(g13782,I16117);
  IV  NOT_5106(g17575,g14921);
  IV  NOT_5107(g28137,I26638);
  IV  NOT_5108(g11984,g9186);
  IV  NOT_5109(g16967,I18125);
  IV  NOT_5110(I22331,g19417);
  IV  NOT_5111(g32668,g31070);
  IV  NOT_5112(g32842,g31710);
  IV  NOT_5113(g17711,I18694);
  IV  NOT_5114(g7046,g5791);
  IV  NOT_5115(I32284,g34052);
  IV  NOT_5116(g20653,I20747);
  IV  NOT_5117(g27991,g25852);
  IV  NOT_5118(I33288,g34989);
  IV  NOT_5119(g31802,g29385);
  IV  NOT_5120(g9631,g6573);
  IV  NOT_5121(g17327,I18310);
  IV  NOT_5122(g25060,g23708);
  IV  NOT_5123(g32489,g30614);
  IV  NOT_5124(g8389,g3125);
  IV  NOT_5125(I13329,g86);
  IV  NOT_5126(I27388,g27698);
  IV  NOT_5127(g31857,g29385);
  IV  NOT_5128(g7446,g1256);
  IV  NOT_5129(g18200,I19012);
  IV  NOT_5130(g29811,g28376);
  IV  NOT_5131(g23223,g21308);
  IV  NOT_5132(g7514,g6704);
  IV  NOT_5133(g19360,g16249);
  IV  NOT_5134(g11418,I14424);
  IV  NOT_5135(g34714,I32874);
  IV  NOT_5136(g8990,g146);
  IV  NOT_5137(g12882,g10389);
  IV  NOT_5138(g9257,g5115);
  IV  NOT_5139(g22492,g19614);
  IV  NOT_5140(g25197,g23958);
  IV  NOT_5141(g29343,g28174);
  IV  NOT_5142(g7003,g5152);
  IV  NOT_5143(I13539,g6381);
  IV  NOT_5144(g22303,g19277);
  IV  NOT_5145(I27777,g29043);
  IV  NOT_5146(g9817,I13374);
  IV  NOT_5147(g32559,g30825);
  IV  NOT_5148(g34315,g34085);
  IV  NOT_5149(g10475,g8844);
  IV  NOT_5150(I17932,g3310);
  IV  NOT_5151(g24138,g21143);
  IV  NOT_5152(g32525,g31170);
  IV  NOT_5153(g32488,g31194);
  IV  NOT_5154(g11170,g8476);
  IV  NOT_5155(g34910,g34864);
  IV  NOT_5156(I29444,g30928);
  IV  NOT_5157(g8171,g3817);
  IV  NOT_5158(g10727,I14016);
  IV  NOT_5159(g7345,g6415);
  IV  NOT_5160(g7841,g904);
  IV  NOT_5161(I12534,g50);
  IV  NOT_5162(g20636,g18008);
  IV  NOT_5163(I19384,g15085);
  IV  NOT_5164(g8787,I12773);
  IV  NOT_5165(g32558,g30735);
  IV  NOT_5166(g34202,I32161);
  IV  NOT_5167(g23084,g19954);
  IV  NOT_5168(g24636,g23121);
  IV  NOT_5169(g6826,g218);
  IV  NOT_5170(g10222,g4492);
  IV  NOT_5171(g7191,g6398);
  IV  NOT_5172(g30055,g29157);
  IV  NOT_5173(g17606,g14999);
  IV  NOT_5174(g20852,g15595);
  IV  NOT_5175(g32830,g31327);
  IV  NOT_5176(g23922,g18997);
  IV  NOT_5177(g23321,I22422);
  IV  NOT_5178(g32893,g30937);
  IV  NOT_5179(I18028,g13638);
  IV  NOT_5180(g21179,g15373);
  IV  NOT_5181(I24920,g25513);
  IV  NOT_5182(g26801,I25511);
  IV  NOT_5183(I24434,g22763);
  IV  NOT_5184(g29368,I27730);
  IV  NOT_5185(g9751,g1710);
  IV  NOT_5186(g34070,g33725);
  IV  NOT_5187(g8281,g3494);
  IV  NOT_5188(g32544,g30735);
  IV  NOT_5189(g19629,g17015);
  IV  NOT_5190(g32865,g31327);
  IV  NOT_5191(g19451,g15938);
  IV  NOT_5192(g21178,g17955);
  IV  NOT_5193(g34590,I32678);
  IV  NOT_5194(g19472,g16349);
  IV  NOT_5195(g24963,g22342);
  IV  NOT_5196(g20664,g15373);
  IV  NOT_5197(g34986,I33258);
  IV  NOT_5198(g32713,g30673);
  IV  NOT_5199(g7536,g5976);
  IV  NOT_5200(g9585,g1616);
  IV  NOT_5201(g8297,g142);
  IV  NOT_5202(g10347,I13759);
  IV  NOT_5203(g21685,I21246);
  IV  NOT_5204(I16733,g12026);
  IV  NOT_5205(I12997,g351);
  IV  NOT_5206(g28726,g27937);
  IV  NOT_5207(g34384,I32391);
  IV  NOT_5208(g23953,g19277);
  IV  NOT_5209(g30067,g29060);
  IV  NOT_5210(g11401,g7593);
  IV  NOT_5211(g22840,g20330);
  IV  NOT_5212(g21654,g17619);
  IV  NOT_5213(I29977,g31596);
  IV  NOT_5214(g7858,g947);
  IV  NOT_5215(g32610,g31070);
  IV  NOT_5216(g20576,g18065);
  IV  NOT_5217(g20585,g17955);
  IV  NOT_5218(g23654,g20248);
  IV  NOT_5219(I12061,g562);
  IV  NOT_5220(g32705,g30614);
  IV  NOT_5221(g34094,g33772);
  IV  NOT_5222(g13477,I15954);
  IV  NOT_5223(g8745,g744);
  IV  NOT_5224(g28436,I26929);
  IV  NOT_5225(g8138,g1500);
  IV  NOT_5226(g8639,g2807);
  IV  NOT_5227(g24585,g23063);
  IV  NOT_5228(I22149,g21036);
  IV  NOT_5229(g19071,g15591);
  IV  NOT_5230(g23800,g21246);
  IV  NOT_5231(I23711,g23192);
  IV  NOT_5232(g20554,g15348);
  IV  NOT_5233(g23417,g20391);
  IV  NOT_5234(g32679,g31579);
  IV  NOT_5235(g16322,I17650);
  IV  NOT_5236(g8791,I12787);
  IV  NOT_5237(g10351,g6802);
  IV  NOT_5238(g23936,g19210);
  IV  NOT_5239(g10372,g6900);
  IV  NOT_5240(I23327,g22647);
  IV  NOT_5241(g25202,g23932);
  IV  NOT_5242(g19776,g17015);
  IV  NOT_5243(g19785,g16987);
  IV  NOT_5244(g34150,I32103);
  IV  NOT_5245(I32963,g34650);
  IV  NOT_5246(g16159,g13584);
  IV  NOT_5247(g22192,g19801);
  IV  NOT_5248(g20609,g15373);
  IV  NOT_5249(g28274,I26799);
  IV  NOT_5250(g15171,I17098);
  IV  NOT_5251(g34877,I33103);
  IV  NOT_5252(g10175,g28);
  IV  NOT_5253(I17723,g13177);
  IV  NOT_5254(g12082,g9645);
  IV  NOT_5255(g17390,g14755);
  IV  NOT_5256(g28593,g27727);
  IV  NOT_5257(g32678,g31528);
  IV  NOT_5258(g13022,g11894);
  IV  NOT_5259(g7522,g6661);
  IV  NOT_5260(g23334,g20785);
  IV  NOT_5261(g25055,g23590);
  IV  NOT_5262(g19147,I19786);
  IV  NOT_5263(g30019,g29060);
  IV  NOT_5264(g7115,g12);
  IV  NOT_5265(g12107,g9687);
  IV  NOT_5266(g8808,g595);
  IV  NOT_5267(g19754,g17062);
  IV  NOT_5268(g7315,g1772);
  IV  NOT_5269(g16158,g13555);
  IV  NOT_5270(g20608,g15171);
  IV  NOT_5271(g25111,g23699);
  IV  NOT_5272(g9669,g5092);
  IV  NOT_5273(g19355,g16027);
  IV  NOT_5274(I12360,g528);
  IV  NOT_5275(g25070,g23590);
  IV  NOT_5276(g32460,g31194);
  IV  NOT_5277(g32686,g31579);
  IV  NOT_5278(I22343,g19371);
  IV  NOT_5279(g24115,g20998);
  IV  NOT_5280(g32939,g31327);
  IV  NOT_5281(I18903,g16872);
  IV  NOT_5282(g30018,g28987);
  IV  NOT_5283(g32383,I29913);
  IV  NOT_5284(g19950,g15885);
  IV  NOT_5285(g14063,g11048);
  IV  NOT_5286(g19370,g15915);
  IV  NOT_5287(I19917,g18088);
  IV  NOT_5288(I14046,g9900);
  IV  NOT_5289(I17148,g14442);
  IV  NOT_5290(g16656,I17852);
  IV  NOT_5291(g9772,I13352);
  IV  NOT_5292(I26638,g27965);
  IV  NOT_5293(g20921,g15426);
  IV  NOT_5294(g12345,g7158);
  IV  NOT_5295(I16476,g10430);
  IV  NOT_5296(g14790,I16855);
  IV  NOT_5297(g20052,g17533);
  IV  NOT_5298(g23964,g19147);
  IV  NOT_5299(I23303,g21669);
  IV  NOT_5300(g32938,g30937);
  IV  NOT_5301(g28034,g26365);
  IV  NOT_5302(g33533,I31361);
  IV  NOT_5303(g29310,g28991);
  IV  NOT_5304(g16680,g13223);
  IV  NOT_5305(g24052,g21193);
  IV  NOT_5306(I17104,g12932);
  IV  NOT_5307(g12940,g11744);
  IV  NOT_5308(g17522,g14927);
  IV  NOT_5309(g21423,g15224);
  IV  NOT_5310(g12399,g9920);
  IV  NOT_5311(g9743,I13321);
  IV  NOT_5312(I16555,g10430);
  IV  NOT_5313(g23423,g20871);
  IV  NOT_5314(g8201,g1894);
  IV  NOT_5315(g9890,g6058);
  IV  NOT_5316(g13305,g11048);
  IV  NOT_5317(g6827,g1277);
  IV  NOT_5318(g14873,I16898);
  IV  NOT_5319(g23216,g20924);
  IV  NOT_5320(g11900,I14708);
  IV  NOT_5321(g19996,g17271);
  IV  NOT_5322(g29379,I27749);
  IV  NOT_5323(g29925,g28820);
  IV  NOT_5324(g13809,I16135);
  IV  NOT_5325(I23381,g23322);
  IV  NOT_5326(I15036,g799);
  IV  NOT_5327(g8449,g3752);
  IV  NOT_5328(g12804,g9927);
  IV  NOT_5329(g9011,g1422);
  IV  NOT_5330(g19367,I19851);
  IV  NOT_5331(g19394,g16326);
  IV  NOT_5332(I12451,g3092);
  IV  NOT_5333(g6846,g2152);
  IV  NOT_5334(g9856,g5343);
  IV  NOT_5335(g8575,g291);
  IV  NOT_5336(g13036,g10981);
  IV  NOT_5337(g32875,g31376);
  IV  NOT_5338(g30917,I28897);
  IV  NOT_5339(I14827,g9686);
  IV  NOT_5340(g11560,g7647);
  IV  NOT_5341(g13101,I15736);
  IV  NOT_5342(g14209,g11415);
  IV  NOT_5343(g7880,g1291);
  IV  NOT_5344(g13177,I15782);
  IV  NOT_5345(g34917,I33143);
  IV  NOT_5346(g8715,g4927);
  IV  NOT_5347(g20674,g15277);
  IV  NOT_5348(g7595,I12067);
  IV  NOT_5349(g23543,g21514);
  IV  NOT_5350(g6803,g496);
  IV  NOT_5351(g16966,g14291);
  IV  NOT_5352(g7537,g311);
  IV  NOT_5353(g24184,I23396);
  IV  NOT_5354(I18845,g6711);
  IV  NOT_5355(I32921,g34650);
  IV  NOT_5356(g16631,g14454);
  IV  NOT_5357(g14208,g11563);
  IV  NOT_5358(I18262,g13857);
  IV  NOT_5359(g29944,g28911);
  IV  NOT_5360(g22904,I22111);
  IV  NOT_5361(g23000,g20453);
  IV  NOT_5362(I26578,g26941);
  IV  NOT_5363(g23908,g20739);
  IV  NOT_5364(g17326,I18307);
  IV  NOT_5365(g32837,g31327);
  IV  NOT_5366(g31856,g29385);
  IV  NOT_5367(I13206,g5448);
  IV  NOT_5368(g8833,g794);
  IV  NOT_5369(g30077,g29057);
  IV  NOT_5370(g9992,g5990);
  IV  NOT_5371(g20732,g15595);
  IV  NOT_5372(g23569,g21611);
  IV  NOT_5373(g25196,g22763);
  IV  NOT_5374(g10542,g7196);
  IV  NOT_5375(I31610,g33149);
  IV  NOT_5376(I23390,g23395);
  IV  NOT_5377(g13064,g11705);
  IV  NOT_5378(g24732,g23042);
  IV  NOT_5379(g14453,I16610);
  IV  NOT_5380(g7017,g128);
  IV  NOT_5381(I30992,g32445);
  IV  NOT_5382(g7243,I11892);
  IV  NOT_5383(g19446,I19917);
  IV  NOT_5384(g34597,I32699);
  IV  NOT_5385(I12776,g4207);
  IV  NOT_5386(I13759,g6754);
  IV  NOT_5387(I18191,g14385);
  IV  NOT_5388(g23568,g21611);
  IV  NOT_5389(I33255,g34975);
  IV  NOT_5390(I33189,g34929);
  IV  NOT_5391(g8584,g3639);
  IV  NOT_5392(g8539,g3454);
  IV  NOT_5393(g23242,g21070);
  IV  NOT_5394(I32973,g34714);
  IV  NOT_5395(I29571,g31783);
  IV  NOT_5396(g34689,I32837);
  IV  NOT_5397(I33270,g34982);
  IV  NOT_5398(g34923,I33161);
  IV  NOT_5399(g9863,g5503);
  IV  NOT_5400(I12355,g46);
  IV  NOT_5401(g16289,g13223);
  IV  NOT_5402(g9480,g559);
  IV  NOT_5403(I17228,g13350);
  IV  NOT_5404(g6994,g4933);
  IV  NOT_5405(g21123,g15615);
  IV  NOT_5406(g18100,I18906);
  IV  NOT_5407(g34688,I32834);
  IV  NOT_5408(g9713,g3618);
  IV  NOT_5409(g10607,g10233);
  IV  NOT_5410(g12833,I15448);
  IV  NOT_5411(g22847,g20283);
  IV  NOT_5412(g16309,I17639);
  IV  NOT_5413(I12950,g4287);
  IV  NOT_5414(g23814,g19074);
  IV  NOT_5415(g10320,g817);
  IV  NOT_5416(g32617,g30825);
  IV  NOT_5417(g28575,g27711);
  IV  NOT_5418(g32470,g31566);
  IV  NOT_5419(g10073,g134);
  IV  NOT_5420(I18832,g13782);
  IV  NOT_5421(I31686,g33164);
  IV  NOT_5422(g7328,g2197);
  IV  NOT_5423(g32915,g31710);
  IV  NOT_5424(g10274,g976);
  IV  NOT_5425(g29765,I28014);
  IV  NOT_5426(g10530,g8922);
  IV  NOT_5427(g7542,I12030);
  IV  NOT_5428(I12858,g4340);
  IV  NOT_5429(g28711,g27886);
  IV  NOT_5430(g13009,I15617);
  IV  NOT_5431(g16308,I17636);
  IV  NOT_5432(g9569,g6227);
  IV  NOT_5433(g13665,g11306);
  IV  NOT_5434(g27004,g26131);
  IV  NOT_5435(g30102,g29157);
  IV  NOT_5436(g8362,g194);
  IV  NOT_5437(I13744,g3518);
  IV  NOT_5438(g31831,g29385);
  IV  NOT_5439(g32201,g31509);
  IV  NOT_5440(g24013,g21611);
  IV  NOT_5441(I33030,g34768);
  IV  NOT_5442(I12151,g604);
  IV  NOT_5443(g10122,I13623);
  IV  NOT_5444(g6816,g933);
  IV  NOT_5445(I12172,g2715);
  IV  NOT_5446(g17183,I18221);
  IV  NOT_5447(g17673,g14723);
  IV  NOT_5448(g17847,I18839);
  IV  NOT_5449(I26430,g26856);
  IV  NOT_5450(g13008,g11855);
  IV  NOT_5451(g15656,I17198);
  IV  NOT_5452(I21483,g18726);
  IV  NOT_5453(g20329,g15277);
  IV  NOT_5454(I33267,g34979);
  IV  NOT_5455(g8052,g1211);
  IV  NOT_5456(I18861,g14307);
  IV  NOT_5457(g21293,I21036);
  IV  NOT_5458(g20207,g17015);
  IV  NOT_5459(g23230,I22327);
  IV  NOT_5460(g15680,I17207);
  IV  NOT_5461(g20539,g15483);
  IV  NOT_5462(g25001,g23666);
  IV  NOT_5463(g17062,I18154);
  IV  NOT_5464(g20005,g17433);
  IV  NOT_5465(g13485,g10476);
  IV  NOT_5466(g20328,g15867);
  IV  NOT_5467(g32595,g30825);
  IV  NOT_5468(g32467,g31194);
  IV  NOT_5469(g32494,g30825);
  IV  NOT_5470(g19902,g17200);
  IV  NOT_5471(g24005,I23149);
  IV  NOT_5472(g17509,I18446);
  IV  NOT_5473(g14034,g11048);
  IV  NOT_5474(g19957,g16540);
  IV  NOT_5475(g16816,I18028);
  IV  NOT_5476(g20538,g15348);
  IV  NOT_5477(g9688,g113);
  IV  NOT_5478(g28606,g27762);
  IV  NOT_5479(g6847,g2283);
  IV  NOT_5480(g13555,g12692);
  IV  NOT_5481(g18882,I19674);
  IV  NOT_5482(g32623,g30735);
  IV  NOT_5483(g18991,g16136);
  IV  NOT_5484(I28897,g30155);
  IV  NOT_5485(g19739,g16931);
  IV  NOT_5486(I25391,g24483);
  IV  NOT_5487(g9976,g2537);
  IV  NOT_5488(g17508,I18443);
  IV  NOT_5489(g29317,I27677);
  IV  NOT_5490(g10153,g2417);
  IV  NOT_5491(g23841,g19074);
  IV  NOT_5492(I22096,g19890);
  IV  NOT_5493(g23992,g19210);
  IV  NOT_5494(g32782,g30735);
  IV  NOT_5495(g23391,g20645);
  IV  NOT_5496(g19146,g15574);
  IV  NOT_5497(g19738,g15992);
  IV  NOT_5498(g33080,I30644);
  IV  NOT_5499(g21510,g15647);
  IV  NOT_5500(g23510,g18833);
  IV  NOT_5501(g10409,g7087);
  IV  NOT_5502(g16752,I17976);
  IV  NOT_5503(I21757,g21308);
  IV  NOT_5504(I33218,g34955);
  IV  NOT_5505(I25579,g25297);
  IV  NOT_5506(g16954,I18104);
  IV  NOT_5507(g29129,g27858);
  IV  NOT_5508(g22213,g19147);
  IV  NOT_5509(g19699,I20116);
  IV  NOT_5510(g8504,g3451);
  IV  NOT_5511(g34511,g34419);
  IV  NOT_5512(g10136,g6113);
  IV  NOT_5513(g16643,I17839);
  IV  NOT_5514(g10408,g7049);
  IV  NOT_5515(g9000,g632);
  IV  NOT_5516(g32822,g30937);
  IV  NOT_5517(g13074,I15702);
  IV  NOT_5518(I24191,g22360);
  IV  NOT_5519(g29128,g27800);
  IV  NOT_5520(g14635,I16741);
  IV  NOT_5521(I12227,g34);
  IV  NOT_5522(g13239,g10632);
  IV  NOT_5523(g19698,g16971);
  IV  NOT_5524(g9326,g6203);
  IV  NOT_5525(I15238,g6351);
  IV  NOT_5526(g12951,I15569);
  IV  NOT_5527(g25157,g22498);
  IV  NOT_5528(g23578,I22725);
  IV  NOT_5529(g8070,g3518);
  IV  NOT_5530(g13594,g11012);
  IV  NOT_5531(I16438,g11165);
  IV  NOT_5532(g23014,g20391);
  IV  NOT_5533(I25586,g25537);
  IV  NOT_5534(g8470,I12605);
  IV  NOT_5535(g20100,I20369);
  IV  NOT_5536(g7512,g5283);
  IV  NOT_5537(g34660,g34473);
  IV  NOT_5538(I30983,g32433);
  IV  NOT_5539(g9760,g2315);
  IV  NOT_5540(g20771,g15171);
  IV  NOT_5541(g22311,g18935);
  IV  NOT_5542(g24100,g20857);
  IV  NOT_5543(g26054,g24804);
  IV  NOT_5544(g7490,g2629);
  IV  NOT_5545(I15382,g9071);
  IV  NOT_5546(I14647,g7717);
  IV  NOT_5547(g25231,g22228);
  IV  NOT_5548(g7166,g4311);
  IV  NOT_5549(g20235,g15277);
  IV  NOT_5550(g19427,g16292);
  IV  NOT_5551(I26130,g26510);
  IV  NOT_5552(g11941,I14761);
  IV  NOT_5553(g19366,g15885);
  IV  NOT_5554(I17857,g3969);
  IV  NOT_5555(g32853,g30673);
  IV  NOT_5556(g24683,g23112);
  IV  NOT_5557(g33736,I31597);
  IV  NOT_5558(g11519,g8481);
  IV  NOT_5559(I14999,g10030);
  IV  NOT_5560(g16195,g13437);
  IV  NOT_5561(g34480,I32535);
  IV  NOT_5562(g16489,I17699);
  IV  NOT_5563(g34916,I33140);
  IV  NOT_5564(g13675,g10556);
  IV  NOT_5565(I20861,g16960);
  IV  NOT_5566(g32589,g31070);
  IV  NOT_5567(g7456,g2495);
  IV  NOT_5568(g15224,I17101);
  IV  NOT_5569(g7148,I11835);
  IV  NOT_5570(g6817,g956);
  IV  NOT_5571(g7649,g1345);
  IV  NOT_5572(g22592,I21930);
  IV  NOT_5573(g22756,g20436);
  IV  NOT_5574(g16525,I17723);
  IV  NOT_5575(g15571,g13211);
  IV  NOT_5576(g26942,I25692);
  IV  NOT_5577(g9924,g5644);
  IV  NOT_5578(g10474,g8841);
  IV  NOT_5579(g32588,g30825);
  IV  NOT_5580(g32524,g31070);
  IV  NOT_5581(g9220,g843);
  IV  NOT_5582(g31843,g29385);
  IV  NOT_5583(g32836,g31021);
  IV  NOT_5584(g33696,I31535);
  IV  NOT_5585(g30076,g29085);
  IV  NOT_5586(g30085,g29082);
  IV  NOT_5587(g7851,g921);
  IV  NOT_5588(I33075,g34843);
  IV  NOT_5589(g9779,g5156);
  IV  NOT_5590(g26655,g25492);
  IV  NOT_5591(g13637,g10556);
  IV  NOT_5592(g20515,g15483);
  IV  NOT_5593(g34307,g34087);
  IV  NOT_5594(g23041,g19882);
  IV  NOT_5595(I20388,g17724);
  IV  NOT_5596(g32477,g31566);
  IV  NOT_5597(I18360,g1426);
  IV  NOT_5598(g21275,g15426);
  IV  NOT_5599(g24515,g22689);
  IV  NOT_5600(I31494,g33283);
  IV  NOT_5601(g24991,g22369);
  IV  NOT_5602(I12120,g632);
  IV  NOT_5603(g10109,g135);
  IV  NOT_5604(g30054,g29134);
  IV  NOT_5605(g21430,g15608);
  IV  NOT_5606(g27163,I25869);
  IV  NOT_5607(g34596,I32696);
  IV  NOT_5608(g8406,g232);
  IV  NOT_5609(g17756,g14858);
  IV  NOT_5610(I27738,g28140);
  IV  NOT_5611(g23430,I22547);
  IV  NOT_5612(g23746,g20902);
  IV  NOT_5613(g23493,g21611);
  IV  NOT_5614(g7964,g3155);
  IV  NOT_5615(g7260,I11908);
  IV  NOT_5616(g8635,g2783);
  IV  NOT_5617(g24407,g22594);
  IV  NOT_5618(g34243,I32228);
  IV  NOT_5619(g29697,g28336);
  IV  NOT_5620(g9977,g2667);
  IV  NOT_5621(g19481,g16349);
  IV  NOT_5622(g10108,g120);
  IV  NOT_5623(I14932,g9901);
  IV  NOT_5624(g29995,g28955);
  IV  NOT_5625(I33037,g34770);
  IV  NOT_5626(g34431,I32464);
  IV  NOT_5627(g12012,g9213);
  IV  NOT_5628(g32118,g31008);
  IV  NOT_5629(g15816,I17314);
  IV  NOT_5630(g8766,g572);
  IV  NOT_5631(g18940,I19719);
  IV  NOT_5632(g8087,g1157);
  IV  NOT_5633(I31782,g33219);
  IV  NOT_5634(g32864,g30937);
  IV  NOT_5635(g23237,g20924);
  IV  NOT_5636(I19734,g17725);
  IV  NOT_5637(g7063,g4831);
  IV  NOT_5638(g10606,g10233);
  IV  NOT_5639(g21340,I21074);
  IV  NOT_5640(g32749,g31021);
  IV  NOT_5641(g32616,g30735);
  IV  NOT_5642(g23340,g21070);
  IV  NOT_5643(g23983,g19210);
  IV  NOT_5644(I22128,g19968);
  IV  NOT_5645(g34773,I32963);
  IV  NOT_5646(g9051,g1426);
  IV  NOT_5647(g23684,I22819);
  IV  NOT_5648(g25480,g22228);
  IV  NOT_5649(g34942,g34928);
  IV  NOT_5650(g32748,g31710);
  IV  NOT_5651(I15577,g10430);
  IV  NOT_5652(g8748,g776);
  IV  NOT_5653(g11215,g8285);
  IV  NOT_5654(g19127,I19775);
  IV  NOT_5655(g9451,g5873);
  IV  NOT_5656(g28326,g27414);
  IV  NOT_5657(I32991,g34759);
  IV  NOT_5658(I14505,g10140);
  IV  NOT_5659(I33155,g34897);
  IV  NOT_5660(g13215,g10909);
  IV  NOT_5661(g26131,I25161);
  IV  NOT_5662(g34156,g33907);
  IV  NOT_5663(g13729,g10951);
  IV  NOT_5664(g25550,g22763);
  IV  NOT_5665(g20441,g17873);
  IV  NOT_5666(g20584,g17873);
  IV  NOT_5667(g32704,g31070);
  IV  NOT_5668(I21047,g17429);
  IV  NOT_5669(g10381,g6957);
  IV  NOT_5670(g28040,g26365);
  IV  NOT_5671(g33708,I31555);
  IV  NOT_5672(I33170,g34890);
  IV  NOT_5673(g19490,g16489);
  IV  NOT_5674(g25287,g22228);
  IV  NOT_5675(g34670,I32794);
  IV  NOT_5676(I29939,g31667);
  IV  NOT_5677(g9999,g6109);
  IV  NOT_5678(I17128,g13835);
  IV  NOT_5679(g23517,g21070);
  IV  NOT_5680(g33258,g32296);
  IV  NOT_5681(g32809,g31327);
  IV  NOT_5682(g32900,g30937);
  IV  NOT_5683(g25307,g22763);
  IV  NOT_5684(g32466,g31070);
  IV  NOT_5685(g7118,g832);
  IV  NOT_5686(g7619,g1296);
  IV  NOT_5687(g16124,g13555);
  IV  NOT_5688(I19487,g15125);
  IV  NOT_5689(g19376,g17509);
  IV  NOT_5690(g19385,g16326);
  IV  NOT_5691(I17626,g14582);
  IV  NOT_5692(g17413,I18350);
  IV  NOT_5693(g9103,g5774);
  IV  NOT_5694(g32808,g30937);
  IV  NOT_5695(I26952,g27972);
  IV  NOT_5696(g24759,g23003);
  IV  NOT_5697(I18071,g13680);
  IV  NOT_5698(g19980,g17226);
  IV  NOT_5699(g25243,g22763);
  IV  NOT_5700(g34839,I33053);
  IV  NOT_5701(g17691,I18674);
  IV  NOT_5702(g20114,I20385);
  IV  NOT_5703(g16686,I17892);
  IV  NOT_5704(g34930,I33182);
  IV  NOT_5705(g11349,I14365);
  IV  NOT_5706(g34993,I33279);
  IV  NOT_5707(g12946,I15564);
  IV  NOT_5708(g15842,g13469);
  IV  NOT_5709(g32560,g31070);
  IV  NOT_5710(g20435,g15348);
  IV  NOT_5711(g8373,g2485);
  IV  NOT_5712(I15906,g10430);
  IV  NOT_5713(g24114,g20720);
  IV  NOT_5714(g8091,g1579);
  IV  NOT_5715(I33167,g34890);
  IV  NOT_5716(g6772,I11629);
  IV  NOT_5717(g29498,I27784);
  IV  NOT_5718(g24082,g19890);
  IV  NOT_5719(I15284,g6697);
  IV  NOT_5720(g16030,g13570);
  IV  NOT_5721(g7393,g5320);
  IV  NOT_5722(g13906,I16201);
  IV  NOT_5723(g10390,g6987);
  IV  NOT_5724(g21362,g17873);
  IV  NOT_5725(g24107,g20857);
  IV  NOT_5726(g32642,g31542);
  IV  NOT_5727(g9732,g5481);
  IV  NOT_5728(g23362,I22467);
  IV  NOT_5729(g34131,I32074);
  IV  NOT_5730(g29056,g27800);
  IV  NOT_5731(g22928,I22131);
  IV  NOT_5732(g9753,g1890);
  IV  NOT_5733(I26516,g26824);
  IV  NOT_5734(g23523,g21514);
  IV  NOT_5735(g31810,g29385);
  IV  NOT_5736(g8283,I12493);
  IV  NOT_5737(g25773,g24453);
  IV  NOT_5738(I27481,g27928);
  IV  NOT_5739(g18833,I19661);
  IV  NOT_5740(g31657,I29239);
  IV  NOT_5741(g7971,g4818);
  IV  NOT_5742(g13304,I15872);
  IV  NOT_5743(I20447,g16244);
  IV  NOT_5744(I28582,g30116);
  IV  NOT_5745(I18825,g6019);
  IV  NOT_5746(I18370,g14873);
  IV  NOT_5747(g24744,g22202);
  IV  NOT_5748(I31477,g33391);
  IV  NOT_5749(g29080,g27779);
  IV  NOT_5750(g7686,g4659);
  IV  NOT_5751(g33375,g32377);
  IV  NOT_5752(g8407,g1171);
  IV  NOT_5753(g17929,I18855);
  IV  NOT_5754(g9072,g2994);
  IV  NOT_5755(g25156,g22498);
  IV  NOT_5756(I29218,g30304);
  IV  NOT_5757(g8920,I12899);
  IV  NOT_5758(g8059,g3171);
  IV  NOT_5759(g32733,g31672);
  IV  NOT_5760(I33119,g34852);
  IV  NOT_5761(g14192,g11385);
  IV  NOT_5762(I18858,g13835);
  IV  NOT_5763(g9472,g6555);
  IV  NOT_5764(g19931,g17200);
  IV  NOT_5765(g25180,g23529);
  IV  NOT_5766(g6856,I11682);
  IV  NOT_5767(I12572,g51);
  IV  NOT_5768(g15830,g13432);
  IV  NOT_5769(g17583,g14968);
  IV  NOT_5770(g8718,g3333);
  IV  NOT_5771(I18151,g13144);
  IV  NOT_5772(g34210,I32173);
  IV  NOT_5773(g32874,g30673);
  IV  NOT_5774(I28925,g29987);
  IV  NOT_5775(g9443,g5489);
  IV  NOT_5776(g21727,I21300);
  IV  NOT_5777(I22512,g19389);
  IV  NOT_5778(g20652,I20744);
  IV  NOT_5779(g28508,I26989);
  IV  NOT_5780(g32630,g30735);
  IV  NOT_5781(g7121,I11820);
  IV  NOT_5782(g23863,g19210);
  IV  NOT_5783(g32693,g31579);
  IV  NOT_5784(I31616,g33219);
  IV  NOT_5785(g21222,g17430);
  IV  NOT_5786(I23396,g23427);
  IV  NOT_5787(g7670,g4104);
  IV  NOT_5788(g23222,g20785);
  IV  NOT_5789(I18367,g13010);
  IV  NOT_5790(g26187,I25190);
  IV  NOT_5791(g29342,g28188);
  IV  NOT_5792(g9316,g5742);
  IV  NOT_5793(g25930,I25028);
  IV  NOT_5794(g7625,I12109);
  IV  NOT_5795(g32665,g31579);
  IV  NOT_5796(I31748,g33228);
  IV  NOT_5797(I13473,g4157);
  IV  NOT_5798(g19520,g16826);
  IV  NOT_5799(g6992,g4899);
  IV  NOT_5800(g12760,g10272);
  IV  NOT_5801(g9434,g5385);
  IV  NOT_5802(g13138,I15765);
  IV  NOT_5803(g17787,I18795);
  IV  NOT_5804(g7232,g4411);
  IV  NOT_5805(g10553,g8971);
  IV  NOT_5806(g25838,g25250);
  IV  NOT_5807(I27784,g29013);
  IV  NOT_5808(I15636,g12075);
  IV  NOT_5809(I33276,g34985);
  IV  NOT_5810(I33285,g34988);
  IV  NOT_5811(g18947,g16136);
  IV  NOT_5812(I27385,g27438);
  IV  NOT_5813(g30039,g29134);
  IV  NOT_5814(g30306,g28796);
  IV  NOT_5815(g25131,g23699);
  IV  NOT_5816(I33053,g34778);
  IV  NOT_5817(g15705,g13217);
  IV  NOT_5818(g26937,I25683);
  IV  NOT_5819(g17302,I18285);
  IV  NOT_5820(g32892,g31021);
  IV  NOT_5821(g23347,I22444);
  IV  NOT_5822(g24135,g20720);
  IV  NOT_5823(g32476,g30673);
  IV  NOT_5824(g32485,g31376);
  IV  NOT_5825(g33459,I30995);
  IV  NOT_5826(I31466,g33318);
  IV  NOT_5827(g7909,g936);
  IV  NOT_5828(g30038,g29097);
  IV  NOT_5829(g23253,g21037);
  IV  NOT_5830(I12103,g572);
  IV  NOT_5831(g11852,I14668);
  IV  NOT_5832(g17743,I18734);
  IV  NOT_5833(g9681,g5798);
  IV  NOT_5834(I22499,g21160);
  IV  NOT_5835(g10040,g2652);
  IV  NOT_5836(I22316,g19361);
  IV  NOT_5837(g32555,g30673);
  IV  NOT_5838(I18446,g13028);
  IV  NOT_5839(g14536,I16651);
  IV  NOT_5840(g19860,g17226);
  IV  NOT_5841(g33458,I30992);
  IV  NOT_5842(g7519,g1157);
  IV  NOT_5843(g24361,g22885);
  IV  NOT_5844(g11963,g9153);
  IV  NOT_5845(g25557,g22763);
  IV  NOT_5846(g32570,g31554);
  IV  NOT_5847(g32712,g30614);
  IV  NOT_5848(g25210,g23802);
  IV  NOT_5849(g32914,g31672);
  IV  NOT_5850(I25351,g24466);
  IV  NOT_5851(g9914,g2533);
  IV  NOT_5852(I20355,g17613);
  IV  NOT_5853(g33918,I31782);
  IV  NOT_5854(g23236,g20785);
  IV  NOT_5855(g20500,g17873);
  IV  NOT_5856(g10621,g7567);
  IV  NOT_5857(g34677,I32815);
  IV  NOT_5858(g29365,g29067);
  IV  NOT_5859(g14252,I16438);
  IV  NOT_5860(I22989,g21175);
  IV  NOT_5861(g13664,g11252);
  IV  NOT_5862(g20049,I20318);
  IV  NOT_5863(g23952,g19277);
  IV  NOT_5864(g23351,g20924);
  IV  NOT_5865(g32907,g30937);
  IV  NOT_5866(I31642,g33204);
  IV  NOT_5867(g33079,I30641);
  IV  NOT_5868(g24049,g20014);
  IV  NOT_5869(I14896,g9820);
  IV  NOT_5870(g29960,g28885);
  IV  NOT_5871(g21175,I20951);
  IV  NOT_5872(g22881,I22096);
  IV  NOT_5873(g23821,g19210);
  IV  NOT_5874(g10564,g9462);
  IV  NOT_5875(g15938,I17401);
  IV  NOT_5876(g16075,g13597);
  IV  NOT_5877(g9413,g1744);
  IV  NOT_5878(g19659,g17062);
  IV  NOT_5879(g14564,I16679);
  IV  NOT_5880(g24048,g19968);
  IV  NOT_5881(I11682,g2756);
  IV  NOT_5882(g11576,g8542);
  IV  NOT_5883(I33064,g34784);
  IV  NOT_5884(I25790,g26424);
  IV  NOT_5885(I17989,g14173);
  IV  NOT_5886(g20004,g17249);
  IV  NOT_5887(g13484,g10981);
  IV  NOT_5888(g32567,g31070);
  IV  NOT_5889(g32594,g30735);
  IV  NOT_5890(g19658,g16987);
  IV  NOT_5891(g23264,g21037);
  IV  NOT_5892(g25286,g22228);
  IV  NOT_5893(g16623,g14127);
  IV  NOT_5894(g10183,g2595);
  IV  NOT_5895(I15609,g12013);
  IV  NOT_5896(g7586,I12056);
  IV  NOT_5897(g23516,g20924);
  IV  NOT_5898(g25039,g22498);
  IV  NOT_5899(I28548,g28147);
  IV  NOT_5900(g10397,g7018);
  IV  NOT_5901(g6976,I11750);
  IV  NOT_5902(g14183,g12381);
  IV  NOT_5903(g14673,I16770);
  IV  NOT_5904(g11609,g7660);
  IV  NOT_5905(g9820,g99);
  IV  NOT_5906(g16782,I18006);
  IV  NOT_5907(g12903,g10411);
  IV  NOT_5908(g20613,g15224);
  IV  NOT_5909(I21787,g19422);
  IV  NOT_5910(I22461,g21225);
  IV  NOT_5911(g31817,g29385);
  IV  NOT_5912(g13312,g11048);
  IV  NOT_5913(I18301,g12976);
  IV  NOT_5914(g32941,g30735);
  IV  NOT_5915(g32382,g31657);
  IV  NOT_5916(g11608,g7659);
  IV  NOT_5917(g19644,g17953);
  IV  NOT_5918(g10509,g10233);
  IV  NOT_5919(I18120,g13350);
  IV  NOT_5920(g32519,g30673);
  IV  NOT_5921(I22031,g21387);
  IV  NOT_5922(I27546,g29041);
  IV  NOT_5923(g32185,I29717);
  IV  NOT_5924(g18421,I19235);
  IV  NOT_5925(g14509,I16626);
  IV  NOT_5926(I15921,g12381);
  IV  NOT_5927(g32675,g31070);
  IV  NOT_5928(g8388,g3010);
  IV  NOT_5929(I23357,g23359);
  IV  NOT_5930(g20273,g17128);
  IV  NOT_5931(g20106,g17328);
  IV  NOT_5932(g12563,g9864);
  IV  NOT_5933(g20605,g17955);
  IV  NOT_5934(g21422,g15373);
  IV  NOT_5935(I26409,g26187);
  IV  NOT_5936(g30217,I28458);
  IV  NOT_5937(g8216,g3092);
  IV  NOT_5938(g10851,I14069);
  IV  NOT_5939(I12089,g744);
  IV  NOT_5940(g10872,g7567);
  IV  NOT_5941(g9601,g4005);
  IV  NOT_5942(g23422,g21611);
  IV  NOT_5943(g32518,g30614);
  IV  NOT_5944(I16328,g878);
  IV  NOT_5945(g24106,g19984);
  IV  NOT_5946(g24605,g23139);
  IV  NOT_5947(I14050,g9963);
  IV  NOT_5948(g29043,I27391);
  IV  NOT_5949(I16538,g10417);
  IV  NOT_5950(g13745,I16102);
  IV  NOT_5951(g32637,g30735);
  IV  NOT_5952(g31656,I29236);
  IV  NOT_5953(I20318,g16920);
  IV  NOT_5954(g17249,I18265);
  IV  NOT_5955(I28002,g28153);
  IV  NOT_5956(g32935,g31672);
  IV  NOT_5957(g24463,g23578);
  IV  NOT_5958(I21769,g19402);
  IV  NOT_5959(I17650,g13271);
  IV  NOT_5960(I28128,g28314);
  IV  NOT_5961(g20033,g16579);
  IV  NOT_5962(g31823,g29385);
  IV  NOT_5963(I32613,g34329);
  IV  NOT_5964(g32883,g30735);
  IV  NOT_5965(g17248,I18262);
  IV  NOT_5966(I30641,g32024);
  IV  NOT_5967(I31555,g33212);
  IV  NOT_5968(I14742,g9534);
  IV  NOT_5969(g19411,g16489);
  IV  NOT_5970(g19527,g16349);
  IV  NOT_5971(g17710,g14764);
  IV  NOT_5972(g24033,g19919);
  IV  NOT_5973(I17198,g13809);
  IV  NOT_5974(g12845,g10358);
  IV  NOT_5975(g27990,g26770);
  IV  NOT_5976(g16853,g13584);
  IV  NOT_5977(I12497,g49);
  IV  NOT_5978(g23542,g21514);
  IV  NOT_5979(g9581,g91);
  IV  NOT_5980(g23021,g20283);
  IV  NOT_5981(g23453,I22576);
  IV  NOT_5982(g10213,g6732);
  IV  NOT_5983(I32947,g34659);
  IV  NOT_5984(g12899,g10407);
  IV  NOT_5985(g21726,I21297);
  IV  NOT_5986(g16589,g14082);
  IV  NOT_5987(g25169,g22763);
  IV  NOT_5988(g29955,g28950);
  IV  NOT_5989(g9060,g3355);
  IV  NOT_5990(I32106,g33653);
  IV  NOT_5991(g23913,g19147);
  IV  NOT_5992(g15915,I17392);
  IV  NOT_5993(g9460,g6154);
  IV  NOT_5994(g24795,g23342);
  IV  NOT_5995(g29970,I28199);
  IV  NOT_5996(g7659,I12141);
  IV  NOT_5997(g12898,g10405);
  IV  NOT_5998(g22647,I21959);
  IV  NOT_5999(g17778,I18778);
  IV  NOT_6000(g16588,g13929);
  IV  NOT_6001(g25168,I24334);
  IV  NOT_6002(g23614,g20248);
  IV  NOT_6003(g25410,g22228);
  IV  NOT_6004(g18829,g15171);
  IV  NOT_6005(I12987,g12);
  IV  NOT_6006(I15732,g6692);
  IV  NOT_6007(g8741,g4821);
  IV  NOT_6008(g10047,g5421);
  IV  NOT_6009(I32812,g34588);
  IV  NOT_6010(g19503,g16349);
  IV  NOT_6011(g29878,g28421);
  IV  NOT_6012(g15277,I17104);
  IV  NOT_6013(g21607,g17873);
  IV  NOT_6014(g22999,g20453);
  IV  NOT_6015(g23607,g21611);
  IV  NOT_6016(g21905,I21486);
  IV  NOT_6017(g14205,g12381);
  IV  NOT_6018(g26654,g25275);
  IV  NOT_6019(g20514,g15348);
  IV  NOT_6020(I25530,g25222);
  IV  NOT_6021(g32501,g30825);
  IV  NOT_6022(g32729,g30937);
  IV  NOT_6023(g18828,g17955);
  IV  NOT_6024(g31631,I29221);
  IV  NOT_6025(g10311,g4633);
  IV  NOT_6026(g23320,I22419);
  IV  NOT_6027(g23905,g21514);
  IV  NOT_6028(g9739,g5752);
  IV  NOT_6029(g32577,g31554);
  IV  NOT_6030(g33631,I31459);
  IV  NOT_6031(I14730,g7717);
  IV  NOT_6032(g18946,g16100);
  IV  NOT_6033(g29171,g27937);
  IV  NOT_6034(g21274,g15373);
  IV  NOT_6035(g14912,I16917);
  IV  NOT_6036(g30321,I28572);
  IV  NOT_6037(g23274,g21070);
  IV  NOT_6038(g20507,g15509);
  IV  NOT_6039(g23530,g20248);
  IV  NOT_6040(g22998,g20391);
  IV  NOT_6041(g27832,I26409);
  IV  NOT_6042(I32234,g34126);
  IV  NOT_6043(g34922,I33158);
  IV  NOT_6044(I24281,g23440);
  IV  NOT_6045(g26936,I25680);
  IV  NOT_6046(g15595,I17173);
  IV  NOT_6047(g32728,g31021);
  IV  NOT_6048(g21346,g17821);
  IV  NOT_6049(g25015,g23662);
  IV  NOT_6050(g6977,I11753);
  IV  NOT_6051(I20957,g16228);
  IV  NOT_6052(g19714,g16821);
  IV  NOT_6053(I13240,g5794);
  IV  NOT_6054(g7275,g1728);
  IV  NOT_6055(g22182,I21766);
  IV  NOT_6056(g29967,g28946);
  IV  NOT_6057(g29994,g29049);
  IV  NOT_6058(g34531,I32594);
  IV  NOT_6059(g9995,g6035);
  IV  NOT_6060(I12644,g3689);
  IV  NOT_6061(I11903,g4414);
  IV  NOT_6062(g23565,g21562);
  IV  NOT_6063(g10072,g9);
  IV  NOT_6064(g32438,g30991);
  IV  NOT_6065(I14690,g9340);
  IV  NOT_6066(g8883,g4709);
  IV  NOT_6067(g7615,I12083);
  IV  NOT_6068(g12440,g9985);
  IV  NOT_6069(g27573,g26667);
  IV  NOT_6070(I20562,g16525);
  IV  NOT_6071(g25556,g22763);
  IV  NOT_6072(g24163,I23333);
  IV  NOT_6073(I33176,g34887);
  IV  NOT_6074(g7174,g6052);
  IV  NOT_6075(g19979,g17226);
  IV  NOT_6076(g16748,I17970);
  IV  NOT_6077(g7374,g2227);
  IV  NOT_6078(g12861,g10367);
  IV  NOT_6079(g17651,g14868);
  IV  NOT_6080(g17672,g14720);
  IV  NOT_6081(g34676,I32812);
  IV  NOT_6082(g8217,g3143);
  IV  NOT_6083(I16515,g12477);
  IV  NOT_6084(I17471,g13394);
  IV  NOT_6085(g9390,g5808);
  IV  NOT_6086(g21292,I21033);
  IV  NOT_6087(g11214,g9602);
  IV  NOT_6088(g32906,g31021);
  IV  NOT_6089(g7985,g3506);
  IV  NOT_6090(g16285,I17612);
  IV  NOT_6091(g8466,g1514);
  IV  NOT_6092(I19762,g15732);
  IV  NOT_6093(g22449,g19597);
  IV  NOT_6094(g34654,I32766);
  IV  NOT_6095(g20541,g17821);
  IV  NOT_6096(I12855,g4311);
  IV  NOT_6097(g16305,g13346);
  IV  NOT_6098(g10350,g6800);
  IV  NOT_6099(g13329,I15893);
  IV  NOT_6100(g16053,I17442);
  IV  NOT_6101(g9501,g5731);
  IV  NOT_6102(g6999,g86);
  IV  NOT_6103(g16809,g14387);
  IV  NOT_6104(g21409,g18008);
  IV  NOT_6105(g22897,g21024);
  IV  NOT_6106(g7239,g5033);
  IV  NOT_6107(I12411,g4809);
  IV  NOT_6108(g23409,g21514);
  IV  NOT_6109(g8165,g3530);
  IV  NOT_6110(g32622,g31376);
  IV  NOT_6111(g8571,g57);
  IV  NOT_6112(g8365,g2060);
  IV  NOT_6113(I26381,g26851);
  IV  NOT_6114(g24789,g23309);
  IV  NOT_6115(g32566,g30825);
  IV  NOT_6116(g19741,g16987);
  IV  NOT_6117(I30537,g32027);
  IV  NOT_6118(g29079,g27742);
  IV  NOT_6119(g7380,g2331);
  IV  NOT_6120(g21408,g15373);
  IV  NOT_6121(g10152,g2122);
  IV  NOT_6122(g7591,g6668);
  IV  NOT_6123(g23408,g21468);
  IV  NOT_6124(g8055,g1236);
  IV  NOT_6125(g10396,g6997);
  IV  NOT_6126(g20325,g15171);
  IV  NOT_6127(g24359,g22550);
  IV  NOT_6128(g19067,g15979);
  IV  NOT_6129(g20920,g15426);
  IV  NOT_6130(g20535,g17847);
  IV  NOT_6131(I13990,g7636);
  IV  NOT_6132(g20434,g18065);
  IV  NOT_6133(g9704,g2575);
  IV  NOT_6134(g31816,g29385);
  IV  NOT_6135(g8133,g4809);
  IV  NOT_6136(g24920,I24089);
  IV  NOT_6137(g24535,g22942);
  IV  NOT_6138(I18376,g14332);
  IV  NOT_6139(g24358,g22550);
  IV  NOT_6140(I18297,g1418);
  IV  NOT_6141(I12503,g215);
  IV  NOT_6142(g17505,g14899);
  IV  NOT_6143(g17404,I18337);
  IV  NOT_6144(g10413,g7110);
  IV  NOT_6145(g8774,g781);
  IV  NOT_6146(g32653,g30825);
  IV  NOT_6147(g19801,I20216);
  IV  NOT_6148(I32473,g34248);
  IV  NOT_6149(g17717,g14937);
  IV  NOT_6150(I17879,g14386);
  IV  NOT_6151(g34423,g34222);
  IV  NOT_6152(g15588,I17166);
  IV  NOT_6153(I22886,g18926);
  IV  NOT_6154(g32138,g31233);
  IV  NOT_6155(I17970,g4027);
  IV  NOT_6156(I20895,g16954);
  IV  NOT_6157(g24121,g20720);
  IV  NOT_6158(I18888,g16644);
  IV  NOT_6159(g8396,g3401);
  IV  NOT_6160(g9250,g1600);
  IV  NOT_6161(g34587,I32671);
  IV  NOT_6162(I13718,g890);
  IV  NOT_6163(g12997,g11826);
  IV  NOT_6164(g10405,g7064);
  IV  NOT_6165(g32636,g31376);
  IV  NOT_6166(I23998,g22182);
  IV  NOT_6167(I32788,g34577);
  IV  NOT_6168(g32415,g31591);
  IV  NOT_6169(g14405,g12170);
  IV  NOT_6170(g19695,g17015);
  IV  NOT_6171(g8538,g3412);
  IV  NOT_6172(I12819,g4277);
  IV  NOT_6173(g29977,g28920);
  IV  NOT_6174(I12910,g4340);
  IV  NOT_6175(g16874,I18066);
  IV  NOT_6176(g32852,g30614);
  IV  NOT_6177(g11235,I14301);
  IV  NOT_6178(I32535,g34296);
  IV  NOT_6179(I25327,g24641);
  IV  NOT_6180(g8509,g4141);
  IV  NOT_6181(g35002,I33300);
  IV  NOT_6182(g19526,g16349);
  IV  NOT_6183(g16630,g14142);
  IV  NOT_6184(g16693,I17901);
  IV  NOT_6185(g26814,g25221);
  IV  NOT_6186(g34543,g34359);
  IV  NOT_6187(I22425,g19379);
  IV  NOT_6188(g24173,I23363);
  IV  NOT_6189(g32963,g30825);
  IV  NOT_6190(g22148,g19074);
  IV  NOT_6191(g7515,I12000);
  IV  NOT_6192(g12871,g10378);
  IV  NOT_6193(g29353,I27713);
  IV  NOT_6194(I12070,g785);
  IV  NOT_6195(I22458,g18954);
  IV  NOT_6196(g23537,g20785);
  IV  NOT_6197(g9568,g6181);
  IV  NOT_6198(g31842,g29385);
  IV  NOT_6199(g32664,g31528);
  IV  NOT_6200(g30569,I28838);
  IV  NOT_6201(I16345,g881);
  IV  NOT_6202(g8418,g2619);
  IV  NOT_6203(I19772,g17818);
  IV  NOT_6204(g34569,I32639);
  IV  NOT_6205(g22646,g19389);
  IV  NOT_6206(I22918,g21451);
  IV  NOT_6207(g17433,I18382);
  IV  NOT_6208(I25606,g25465);
  IV  NOT_6209(g8290,g218);
  IV  NOT_6210(I17425,g13416);
  IV  NOT_6211(g18903,g15758);
  IV  NOT_6212(g30568,g29339);
  IV  NOT_6213(g23283,g20785);
  IV  NOT_6214(g19866,g16540);
  IV  NOT_6215(g11991,g9485);
  IV  NOT_6216(I17919,g14609);
  IV  NOT_6217(g13414,g11048);
  IV  NOT_6218(I22444,g19626);
  IV  NOT_6219(g23492,g21562);
  IV  NOT_6220(g25423,I24558);
  IV  NOT_6221(g23303,g20785);
  IV  NOT_6222(I31622,g33204);
  IV  NOT_6223(g32576,g30614);
  IV  NOT_6224(g24134,g19984);
  IV  NOT_6225(g8093,g1624);
  IV  NOT_6226(g32484,g31566);
  IV  NOT_6227(g34242,I32225);
  IV  NOT_6228(g24029,g20982);
  IV  NOT_6229(g33424,g32415);
  IV  NOT_6230(I11701,g4164);
  IV  NOT_6231(g10113,g2084);
  IV  NOT_6232(g17811,g12925);
  IV  NOT_6233(g17646,I18609);
  IV  NOT_6234(I11777,g5357);
  IV  NOT_6235(g20506,g15426);
  IV  NOT_6236(I28199,g28803);
  IV  NOT_6237(I25750,g26823);
  IV  NOT_6238(g20028,g15371);
  IV  NOT_6239(I12067,g739);
  IV  NOT_6240(I32173,g33645);
  IV  NOT_6241(g32554,g30614);
  IV  NOT_6242(I18089,g13144);
  IV  NOT_6243(g24506,I23711);
  IV  NOT_6244(I20385,g16194);
  IV  NOT_6245(g7750,g1070);
  IV  NOT_6246(g24028,g20841);
  IV  NOT_6247(I24784,g24265);
  IV  NOT_6248(g34123,I32062);
  IV  NOT_6249(g16712,g13223);
  IV  NOT_6250(g26841,g24893);
  IV  NOT_6251(g32609,g30735);
  IV  NOT_6252(g21381,g18008);
  IV  NOT_6253(I27735,g28779);
  IV  NOT_6254(I29239,g29498);
  IV  NOT_6255(g31830,g29385);
  IV  NOT_6256(g23982,g19147);
  IV  NOT_6257(g10357,g6825);
  IV  NOT_6258(g26510,I25369);
  IV  NOT_6259(g14357,g12181);
  IV  NOT_6260(g34772,I32960);
  IV  NOT_6261(I12735,g4572);
  IV  NOT_6262(g8181,g424);
  IV  NOT_6263(g28779,I27253);
  IV  NOT_6264(g32608,g31376);
  IV  NOT_6265(g8381,g2610);
  IV  NOT_6266(g19689,g16795);
  IV  NOT_6267(g7040,g4821);
  IV  NOT_6268(g25117,g22417);
  IV  NOT_6269(I16135,g10430);
  IV  NOT_6270(g25000,g23630);
  IV  NOT_6271(g8685,g1430);
  IV  NOT_6272(g7440,g329);
  IV  NOT_6273(g8700,g4054);
  IV  NOT_6274(g28081,I26584);
  IV  NOT_6275(g32921,g31672);
  IV  NOT_6276(g33713,I31564);
  IV  NOT_6277(g8397,g3470);
  IV  NOT_6278(g19688,g16777);
  IV  NOT_6279(g9626,g6466);
  IV  NOT_6280(g8021,g3512);
  IV  NOT_6281(g16594,I17772);
  IV  NOT_6282(g26835,I25555);
  IV  NOT_6283(g13584,g12735);
  IV  NOT_6284(g18990,g16136);
  IV  NOT_6285(g32745,g31376);
  IV  NOT_6286(I29185,g30012);
  IV  NOT_6287(g22896,g21012);
  IV  NOT_6288(I18700,g6027);
  IV  NOT_6289(g23840,g19074);
  IV  NOT_6290(g15733,I17249);
  IV  NOT_6291(g32799,g31710);
  IV  NOT_6292(g18898,g15566);
  IV  NOT_6293(g23390,g21468);
  IV  NOT_6294(g32813,g31710);
  IV  NOT_6295(g22228,I21810);
  IV  NOT_6296(g6820,g1070);
  IV  NOT_6297(g33705,I31550);
  IV  NOT_6298(g25242,g23684);
  IV  NOT_6299(g7666,g4076);
  IV  NOT_6300(I17159,g13350);
  IV  NOT_6301(g20649,g18065);
  IV  NOT_6302(I17125,g13809);
  IV  NOT_6303(I22561,g20841);
  IV  NOT_6304(I23149,g19061);
  IV  NOT_6305(g31189,I29002);
  IV  NOT_6306(g34992,I33276);
  IV  NOT_6307(I17901,g3976);
  IV  NOT_6308(g34391,g34200);
  IV  NOT_6309(g32798,g31672);
  IV  NOT_6310(I22353,g19375);
  IV  NOT_6311(g28380,g27064);
  IV  NOT_6312(g20240,g17847);
  IV  NOT_6313(I23387,g23394);
  IV  NOT_6314(g32973,g31021);
  IV  NOT_6315(I30904,g32424);
  IV  NOT_6316(g34510,g34418);
  IV  NOT_6317(g22716,g19795);
  IV  NOT_6318(g23192,g20248);
  IV  NOT_6319(g16675,I17873);
  IV  NOT_6320(g20648,g15615);
  IV  NOT_6321(g10881,g7567);
  IV  NOT_6322(I17783,g13304);
  IV  NOT_6323(g20903,g17249);
  IV  NOT_6324(g32805,g31672);
  IV  NOT_6325(g13082,g10981);
  IV  NOT_6326(g32674,g30735);
  IV  NOT_6327(g24648,g23148);
  IV  NOT_6328(g7528,g930);
  IV  NOT_6329(g12859,g10366);
  IV  NOT_6330(g13107,g10476);
  IV  NOT_6331(g34579,I32659);
  IV  NOT_6332(g7648,I12135);
  IV  NOT_6333(g26615,g25432);
  IV  NOT_6334(g12950,g12708);
  IV  NOT_6335(g20604,g17873);
  IV  NOT_6336(g9683,g6140);
  IV  NOT_6337(g23522,g21514);
  IV  NOT_6338(g18832,g15634);
  IV  NOT_6339(I13360,g5343);
  IV  NOT_6340(g24604,g23112);
  IV  NOT_6341(g30578,g29956);
  IV  NOT_6342(g33460,I30998);
  IV  NOT_6343(g33686,g33187);
  IV  NOT_6344(g19885,g17249);
  IV  NOT_6345(g26720,g25275);
  IV  NOT_6346(g7655,g4332);
  IV  NOT_6347(g11744,I14602);
  IV  NOT_6348(g20770,g17955);
  IV  NOT_6349(I26508,g26814);
  IV  NOT_6350(g9778,g5069);
  IV  NOT_6351(I14271,g8456);
  IV  NOT_6352(g20563,g15171);
  IV  NOT_6353(g27996,I26508);
  IV  NOT_6354(g32732,g30825);
  IV  NOT_6355(g24770,g22763);
  IV  NOT_6356(g8631,g283);
  IV  NOT_6357(g25230,g23314);
  IV  NOT_6358(g32934,g30735);
  IV  NOT_6359(g24981,g22763);
  IV  NOT_6360(I24089,g22409);
  IV  NOT_6361(g11849,g7601);
  IV  NOT_6362(I16613,g10430);
  IV  NOT_6363(g17582,g14768);
  IV  NOT_6364(g12996,g11823);
  IV  NOT_6365(g10027,g6523);
  IV  NOT_6366(g23483,g18833);
  IV  NOT_6367(I18060,g14198);
  IV  NOT_6368(I23369,g23347);
  IV  NOT_6369(g14662,I16762);
  IV  NOT_6370(g8301,g1399);
  IV  NOT_6371(g19763,g16431);
  IV  NOT_6372(g25265,I24455);
  IV  NOT_6373(I32240,g34131);
  IV  NOT_6374(g29976,g29018);
  IV  NOT_6375(g12844,g10360);
  IV  NOT_6376(g7410,g2008);
  IV  NOT_6377(g11398,I14409);
  IV  NOT_6378(g23862,g19147);
  IV  NOT_6379(g12367,I15205);
  IV  NOT_6380(g32692,g31528);
  IV  NOT_6381(g32761,g30825);
  IV  NOT_6382(I32648,g34371);
  IV  NOT_6383(g18926,I19707);
  IV  NOT_6384(I18855,g13745);
  IV  NOT_6385(I11629,g19);
  IV  NOT_6386(g11652,g7674);
  IV  NOT_6387(g9661,g3661);
  IV  NOT_6388(g13141,g11374);
  IV  NOT_6389(g29374,I27742);
  IV  NOT_6390(g20767,g17873);
  IV  NOT_6391(g26340,g24953);
  IV  NOT_6392(g21326,I21058);
  IV  NOT_6393(g18099,I18903);
  IV  NOT_6394(I18411,g13018);
  IV  NOT_6395(g30116,I28349);
  IV  NOT_6396(I14650,g9340);
  IV  NOT_6397(g33875,I31727);
  IV  NOT_6398(I24497,g22592);
  IV  NOT_6399(g10710,I14006);
  IV  NOT_6400(g20899,I20861);
  IV  NOT_6401(I12300,g1157);
  IV  NOT_6402(g10003,I13539);
  IV  NOT_6403(g23948,g21012);
  IV  NOT_6404(I32770,g34505);
  IV  NOT_6405(g18098,I18900);
  IV  NOT_6406(g10204,g2685);
  IV  NOT_6407(I29438,g30610);
  IV  NOT_6408(g21904,I21483);
  IV  NOT_6409(g14204,g12155);
  IV  NOT_6410(g16577,I17747);
  IV  NOT_6411(g20633,g15171);
  IV  NOT_6412(g23904,g18997);
  IV  NOT_6413(I16371,g887);
  IV  NOT_6414(g31837,g29385);
  IV  NOT_6415(g14779,I16847);
  IV  NOT_6416(g21252,g15656);
  IV  NOT_6417(I22289,g19446);
  IV  NOT_6418(g32329,g31522);
  IV  NOT_6419(g29669,I27941);
  IV  NOT_6420(g34275,g34047);
  IV  NOT_6421(g19480,g16349);
  IV  NOT_6422(g23252,I22353);
  IV  NOT_6423(g17603,g14993);
  IV  NOT_6424(g20191,g17821);
  IV  NOT_6425(g34430,I32461);
  IV  NOT_6426(g17742,g14971);
  IV  NOT_6427(g32539,g31170);
  IV  NOT_6428(g10081,g2279);
  IV  NOT_6429(g17096,I18168);
  IV  NOT_6430(I18894,g16708);
  IV  NOT_6431(g6995,g4944);
  IV  NOT_6432(g7618,I12092);
  IV  NOT_6433(g8441,g3361);
  IV  NOT_6434(g22857,g20739);
  IV  NOT_6435(I22571,g20097);
  IV  NOT_6436(I11785,g5703);
  IV  NOT_6437(g7235,g4521);
  IV  NOT_6438(g7343,g5290);
  IV  NOT_6439(I14365,g3303);
  IV  NOT_6440(g30237,I28480);
  IV  NOT_6441(I16795,g5637);
  IV  NOT_6442(g25007,g22457);
  IV  NOT_6443(g32538,g31070);
  IV  NOT_6444(g24718,g22182);
  IV  NOT_6445(I32794,g34580);
  IV  NOT_6446(g14786,g12471);
  IV  NOT_6447(g29195,I27495);
  IV  NOT_6448(g9484,g1612);
  IV  NOT_6449(g30983,g29657);
  IV  NOT_6450(g9439,g5428);
  IV  NOT_6451(g17681,g14735);
  IV  NOT_6452(g7566,I12049);
  IV  NOT_6453(g6840,g1992);
  IV  NOT_6454(g8673,g4737);
  IV  NOT_6455(g16349,I17661);
  IV  NOT_6456(g34983,I33249);
  IV  NOT_6457(g18997,I19756);
  IV  NOT_6458(g10356,g6819);
  IV  NOT_6459(g33455,I30983);
  IV  NOT_6460(g21183,g15509);
  IV  NOT_6461(g21673,I21234);
  IV  NOT_6462(g7693,g4849);
  IV  NOT_6463(g11833,g8026);
  IV  NOT_6464(g17429,I18370);
  IV  NOT_6465(g7134,g5029);
  IV  NOT_6466(g21397,g15171);
  IV  NOT_6467(g23847,g19210);
  IV  NOT_6468(g13049,I15677);
  IV  NOT_6469(g10380,g6960);
  IV  NOT_6470(g30142,g28754);
  IV  NOT_6471(g18061,g14800);
  IV  NOT_6472(g16284,I17609);
  IV  NOT_6473(g19431,g16249);
  IV  NOT_6474(g34142,I32089);
  IV  NOT_6475(g25116,g22369);
  IV  NOT_6476(g17428,I18367);
  IV  NOT_6477(I22816,g19862);
  IV  NOT_6478(g7548,g1036);
  IV  NOT_6479(g11048,I14158);
  IV  NOT_6480(g8669,g3767);
  IV  NOT_6481(g10090,g5348);
  IV  NOT_6482(g20573,g17384);
  IV  NOT_6483(g10233,I13699);
  IV  NOT_6484(g20247,g17015);
  IV  NOT_6485(g29893,g28755);
  IV  NOT_6486(I24060,g22202);
  IV  NOT_6487(g16622,g14104);
  IV  NOT_6488(g23509,g21611);
  IV  NOT_6489(g10182,g2681);
  IV  NOT_6490(g28620,g27679);
  IV  NOT_6491(I21959,g20242);
  IV  NOT_6492(g20389,g15277);
  IV  NOT_6493(g8058,g3115);
  IV  NOT_6494(I14708,g9417);
  IV  NOT_6495(I28458,g28443);
  IV  NOT_6496(I29139,g29382);
  IV  NOT_6497(g8531,g3288);
  IV  NOT_6498(g19773,g17615);
  IV  NOT_6499(g24389,g22908);
  IV  NOT_6500(g8458,g294);
  IV  NOT_6501(g24045,g21193);
  IV  NOT_6502(g12902,g10409);
  IV  NOT_6503(g20612,g18008);
  IV  NOT_6504(g23508,g21562);
  IV  NOT_6505(I16163,g11930);
  IV  NOT_6506(I20870,g16216);
  IV  NOT_6507(g32771,g31021);
  IV  NOT_6508(g8743,g550);
  IV  NOT_6509(g20388,g17297);
  IV  NOT_6510(g20324,g17955);
  IV  NOT_6511(g8890,g376);
  IV  NOT_6512(I23378,g23426);
  IV  NOT_6513(g29713,I27970);
  IV  NOT_6514(g24099,g20720);
  IV  NOT_6515(g24388,g22885);
  IV  NOT_6516(g20701,g17955);
  IV  NOT_6517(g20777,g15224);
  IV  NOT_6518(g20534,g17183);
  IV  NOT_6519(g22317,g19801);
  IV  NOT_6520(g31623,g29669);
  IV  NOT_6521(g32683,g30614);
  IV  NOT_6522(I17976,g13638);
  IV  NOT_6523(g25465,g23824);
  IV  NOT_6524(g19670,g16897);
  IV  NOT_6525(g24534,g22670);
  IV  NOT_6526(g8505,g3480);
  IV  NOT_6527(g20272,g17239);
  IV  NOT_6528(g34130,I32071);
  IV  NOT_6529(g24098,g19984);
  IV  NOT_6530(g14331,I16489);
  IV  NOT_6531(g12738,g9374);
  IV  NOT_6532(I19863,g16675);
  IV  NOT_6533(g9616,g5452);
  IV  NOT_6534(g17504,g15021);
  IV  NOT_6535(I16541,g11929);
  IV  NOT_6536(g8011,g3167);
  IV  NOT_6537(g25340,g22763);
  IV  NOT_6538(g25035,g23699);
  IV  NOT_6539(I17374,g13638);
  IV  NOT_6540(g8411,I12577);
  IV  NOT_6541(g8734,g4045);
  IV  NOT_6542(g19734,g16861);
  IV  NOT_6543(g13106,g10981);
  IV  NOT_6544(g27698,g26648);
  IV  NOT_6545(g29042,I27388);
  IV  NOT_6546(g13605,I16040);
  IV  NOT_6547(g10897,g7601);
  IV  NOT_6548(I33214,g34954);
  IV  NOT_6549(I20867,g16216);
  IV  NOT_6550(I27314,g28009);
  IV  NOT_6551(g6954,g4138);
  IV  NOT_6552(g19930,g17200);
  IV  NOT_6553(g6810,g723);
  IV  NOT_6554(g9527,g6500);
  IV  NOT_6555(I14069,g9104);
  IV  NOT_6556(g11812,g7567);
  IV  NOT_6557(g7202,g4639);
  IV  NOT_6558(I16724,g12108);
  IV  NOT_6559(g10404,g7026);
  IV  NOT_6560(I12314,g1500);
  IV  NOT_6561(g13463,g10476);
  IV  NOT_6562(g31822,g29385);
  IV  NOT_6563(g32515,g30825);
  IV  NOT_6564(I31539,g33212);
  IV  NOT_6565(g32882,g31376);
  IV  NOT_6566(I14602,g9340);
  IV  NOT_6567(I15033,g10273);
  IV  NOT_6568(g19694,g16429);
  IV  NOT_6569(g7908,g4157);
  IV  NOT_6570(I32388,g34153);
  IV  NOT_6571(g24032,g21256);
  IV  NOT_6572(g22626,I21941);
  IV  NOT_6573(I21802,g21308);
  IV  NOT_6574(I16829,g6715);
  IV  NOT_6575(g25517,g22228);
  IV  NOT_6576(g11033,g8500);
  IV  NOT_6577(g11371,g7565);
  IV  NOT_6578(I16535,g11235);
  IV  NOT_6579(g18911,g15169);
  IV  NOT_6580(g23452,g21468);
  IV  NOT_6581(g10026,g6494);
  IV  NOT_6582(g32407,I29939);
  IV  NOT_6583(g9546,g2437);
  IV  NOT_6584(g13033,g11917);
  IV  NOT_6585(g21205,g15656);
  IV  NOT_6586(g11234,g8355);
  IV  NOT_6587(g10212,g6390);
  IV  NOT_6588(I14970,g9965);
  IV  NOT_6589(g29939,g28857);
  IV  NOT_6590(g17128,I18180);
  IV  NOT_6591(g7518,g1024);
  IV  NOT_6592(I17668,g13279);
  IV  NOT_6593(I20819,g17088);
  IV  NOT_6594(I22525,g19345);
  IV  NOT_6595(I22488,g18984);
  IV  NOT_6596(I17842,g13051);
  IV  NOT_6597(I20910,g17197);
  IV  NOT_6598(g16963,I18117);
  IV  NOT_6599(g23912,g19147);
  IV  NOT_6600(I17392,g13680);
  IV  NOT_6601(g34222,I32195);
  IV  NOT_6602(g9970,g1714);
  IV  NOT_6603(g24061,g19919);
  IV  NOT_6604(I29585,g31655);
  IV  NOT_6605(g29093,g27858);
  IV  NOT_6606(g34437,I32482);
  IV  NOT_6607(g20766,g17433);
  IV  NOT_6608(I26929,g27980);
  IV  NOT_6609(g8080,g3863);
  IV  NOT_6610(I18526,g13055);
  IV  NOT_6611(g31853,g29385);
  IV  NOT_6612(g19502,g15674);
  IV  NOT_6613(g8480,g3147);
  IV  NOT_6614(g19210,I19796);
  IV  NOT_6615(g17533,I18482);
  IV  NOT_6616(g25193,g22763);
  IV  NOT_6617(g8713,g4826);
  IV  NOT_6618(g21051,g15171);
  IV  NOT_6619(g7593,I12061);
  IV  NOT_6620(I17488,g13394);
  IV  NOT_6621(g15348,I17111);
  IV  NOT_6622(g19618,g16349);
  IV  NOT_6623(g19443,g16449);
  IV  NOT_6624(I14967,g9964);
  IV  NOT_6625(g12895,g10403);
  IV  NOT_6626(I12773,g4204);
  IV  NOT_6627(g16585,g14075);
  IV  NOT_6628(g13514,I15987);
  IV  NOT_6629(g25523,g22550);
  IV  NOT_6630(g31836,g29385);
  IV  NOT_6631(g32441,I29969);
  IV  NOT_6632(g32584,g30673);
  IV  NOT_6633(I32997,g34760);
  IV  NOT_6634(g24360,g22228);
  IV  NOT_6635(g29219,I27573);
  IV  NOT_6636(g15566,I17143);
  IV  NOT_6637(g20447,g15426);
  IV  NOT_6638(g14149,g12381);
  IV  NOT_6639(g10387,g6996);
  IV  NOT_6640(g16609,g14454);
  IV  NOT_6641(g19469,g16326);
  IV  NOT_6642(I28336,g29147);
  IV  NOT_6643(g10620,g10233);
  IV  NOT_6644(g17737,g14810);
  IV  NOT_6645(g22856,g20453);
  IV  NOT_6646(g29218,I27570);
  IV  NOT_6647(g22995,g20330);
  IV  NOT_6648(g32759,g31376);
  IV  NOT_6649(g16200,g13584);
  IV  NOT_6650(I33235,g34957);
  IV  NOT_6651(g23350,g20785);
  IV  NOT_6652(g25006,g22417);
  IV  NOT_6653(g32725,g30825);
  IV  NOT_6654(g24162,I23330);
  IV  NOT_6655(I32766,g34522);
  IV  NOT_6656(g7933,g907);
  IV  NOT_6657(g16608,g14116);
  IV  NOT_6658(g19468,g15938);
  IV  NOT_6659(g9617,I13240);
  IV  NOT_6660(g23820,g19147);
  IV  NOT_6661(g34952,g34942);
  IV  NOT_6662(g34351,g34174);
  IV  NOT_6663(g13012,I15626);
  IV  NOT_6664(g32758,g31327);
  IV  NOT_6665(g7521,g5630);
  IV  NOT_6666(I32871,g34521);
  IV  NOT_6667(g25222,I24400);
  IV  NOT_6668(g7050,g5845);
  IV  NOT_6669(g20629,g17955);
  IV  NOT_6670(g23152,g20283);
  IV  NOT_6671(I12930,g4349);
  IV  NOT_6672(I13699,g4581);
  IV  NOT_6673(g9516,g6116);
  IV  NOT_6674(I21002,g16709);
  IV  NOT_6675(g20451,g15277);
  IV  NOT_6676(g21396,g17955);
  IV  NOT_6677(g31616,I29214);
  IV  NOT_6678(I14079,g7231);
  IV  NOT_6679(g30063,g29015);
  IV  NOT_6680(I22124,g21300);
  IV  NOT_6681(g9771,g3969);
  IV  NOT_6682(I29973,g31213);
  IV  NOT_6683(g26834,I25552);
  IV  NOT_6684(g20911,g15171);
  IV  NOT_6685(I16028,g12381);
  IV  NOT_6686(g10369,g6873);
  IV  NOT_6687(g32744,g31327);
  IV  NOT_6688(I31515,g33187);
  IV  NOT_6689(g24911,I24078);
  IV  NOT_6690(g19677,g17096);
  IV  NOT_6691(I18280,g12951);
  IV  NOT_6692(g12490,I15316);
  IV  NOT_6693(g17512,g12983);
  IV  NOT_6694(I17679,g13416);
  IV  NOT_6695(g21413,g15585);
  IV  NOT_6696(g9299,g5124);
  IV  NOT_6697(I15788,g10430);
  IV  NOT_6698(g23413,g21012);
  IV  NOT_6699(g27956,I26466);
  IV  NOT_6700(g32849,g31021);
  IV  NOT_6701(g9547,g2735);
  IV  NOT_6702(g10368,g6887);
  IV  NOT_6703(g32940,g31376);
  IV  NOT_6704(g7379,g2299);
  IV  NOT_6705(g8400,g4836);
  IV  NOT_6706(g11724,I14593);
  IV  NOT_6707(I17188,g13782);
  IV  NOT_6708(g31809,g29385);
  IV  NOT_6709(I12487,g3443);
  IV  NOT_6710(g11325,g7543);
  IV  NOT_6711(g20071,g16826);
  IV  NOT_6712(g32848,g30825);
  IV  NOT_6713(g9892,g6428);
  IV  NOT_6714(g24071,g20841);
  IV  NOT_6715(g11829,I14653);
  IV  NOT_6716(g12889,g10396);
  IV  NOT_6717(g11920,I14730);
  IV  NOT_6718(I11632,g16);
  IV  NOT_6719(g20591,g15509);
  IV  NOT_6720(g25781,g24510);
  IV  NOT_6721(g10412,g7072);
  IV  NOT_6722(g20776,g18008);
  IV  NOT_6723(g20785,I20846);
  IV  NOT_6724(g31808,g29385);
  IV  NOT_6725(g32652,g30735);
  IV  NOT_6726(g32804,g30735);
  IV  NOT_6727(g14412,I16564);
  IV  NOT_6728(g7289,g4382);
  IV  NOT_6729(I12618,g3338);
  IV  NOT_6730(g12888,g10395);
  IV  NOT_6731(g26614,g25426);
  IV  NOT_6732(g10133,g6049);
  IV  NOT_6733(g20147,g17328);
  IV  NOT_6734(I17938,g3676);
  IV  NOT_6735(g34209,I32170);
  IV  NOT_6736(g7835,g4125);
  IV  NOT_6737(g24147,g19402);
  IV  NOT_6738(g10229,g6736);
  IV  NOT_6739(I18066,g3317);
  IV  NOT_6740(g12181,g9478);
  IV  NOT_6741(g26607,g25382);
  IV  NOT_6742(g17499,g14885);
  IV  NOT_6743(g22989,g20453);
  IV  NOT_6744(g23929,g19147);
  IV  NOT_6745(g17316,I18293);
  IV  NOT_6746(g11344,g9015);
  IV  NOT_6747(g34208,g33838);
  IV  NOT_6748(I14158,g8806);
  IV  NOT_6749(g19410,g16449);
  IV  NOT_6750(g24825,g23204);
  IV  NOT_6751(g22722,I22031);
  IV  NOT_6752(g17498,g14688);
  IV  NOT_6753(g22988,g20391);
  IV  NOT_6754(g8183,g482);
  IV  NOT_6755(g23020,g19869);
  IV  NOT_6756(I15682,g12182);
  IV  NOT_6757(g23928,g21562);
  IV  NOT_6758(g8608,g278);
  IV  NOT_6759(I18885,g16643);
  IV  NOT_6760(g30021,g28994);
  IV  NOT_6761(I32071,g33665);
  IV  NOT_6762(g19479,g16449);
  IV  NOT_6763(g19666,g17188);
  IV  NOT_6764(g6782,I11632);
  IV  NOT_6765(g25264,g23828);
  IV  NOT_6766(g16692,g14170);
  IV  NOT_6767(g25790,g25027);
  IV  NOT_6768(I29013,g29705);
  IV  NOT_6769(g25137,g22432);
  IV  NOT_6770(g9340,I13094);
  IV  NOT_6771(I13715,g71);
  IV  NOT_6772(g17056,g13437);
  IV  NOT_6773(I29214,g30300);
  IV  NOT_6774(g11291,g7526);
  IV  NOT_6775(I32591,g34287);
  IV  NOT_6776(g24172,I23360);
  IV  NOT_6777(g23046,g20283);
  IV  NOT_6778(g32962,g30735);
  IV  NOT_6779(g9478,I13152);
  IV  NOT_6780(I14823,g8056);
  IV  NOT_6781(g19478,g16000);
  IV  NOT_6782(g24996,g22763);
  IV  NOT_6783(g17611,g14822);
  IV  NOT_6784(g17722,I18709);
  IV  NOT_6785(g9907,g1959);
  IV  NOT_6786(g13173,g10632);
  IV  NOT_6787(g34913,I33131);
  IV  NOT_6788(g10582,g7116);
  IV  NOT_6789(I16755,g12377);
  IV  NOT_6790(I29207,g30293);
  IV  NOT_6791(g14582,I16698);
  IV  NOT_6792(g33874,I31724);
  IV  NOT_6793(g9959,g6177);
  IV  NOT_6794(g7674,I12151);
  IV  NOT_6795(g8977,g4349);
  IV  NOT_6796(g24367,g22550);
  IV  NOT_6797(g24394,g22228);
  IV  NOT_6798(I16770,g6023);
  IV  NOT_6799(g32500,g30735);
  IV  NOT_6800(g34436,I32479);
  IV  NOT_6801(g9517,g6163);
  IV  NOT_6802(g9690,g732);
  IV  NOT_6803(g17432,I18379);
  IV  NOT_6804(g23787,g18997);
  IV  NOT_6805(I27677,g28156);
  IV  NOT_6806(g29170,g27907);
  IV  NOT_6807(g32833,g30825);
  IV  NOT_6808(g18957,I19734);
  IV  NOT_6809(g21282,I21019);
  IV  NOT_6810(g16214,g13437);
  IV  NOT_6811(g17271,I18270);
  IV  NOT_6812(I32950,g34713);
  IV  NOT_6813(g23282,g20330);
  IV  NOT_6814(I26710,g27511);
  IV  NOT_6815(g7541,g344);
  IV  NOT_6816(g10627,I13968);
  IV  NOT_6817(I25105,g25284);
  IV  NOT_6818(g34320,g34119);
  IV  NOT_6819(g27089,g26703);
  IV  NOT_6820(g10379,g6953);
  IV  NOT_6821(g23302,g20330);
  IV  NOT_6822(I25743,g25903);
  IV  NOT_6823(g31665,I29245);
  IV  NOT_6824(g25209,g22763);
  IV  NOT_6825(g19580,g16164);
  IV  NOT_6826(g30593,g29970);
  IV  NOT_6827(g33665,I31500);
  IV  NOT_6828(g6998,g4932);
  IV  NOT_6829(g22199,g19210);
  IV  NOT_6830(g34530,I32591);
  IV  NOT_6831(g10112,g1988);
  IV  NOT_6832(g34593,I32687);
  IV  NOT_6833(g7132,g4558);
  IV  NOT_6834(g12546,g8740);
  IV  NOT_6835(I22470,g21326);
  IV  NOT_6836(g10050,g6336);
  IV  NOT_6837(g27088,g26694);
  IV  NOT_6838(g18562,I19384);
  IV  NOT_6839(g34346,g34162);
  IV  NOT_6840(g10378,g6926);
  IV  NOT_6841(g25208,g22763);
  IV  NOT_6842(g30565,I28832);
  IV  NOT_6843(g7153,g5373);
  IV  NOT_6844(g7680,g4108);
  IV  NOT_6845(g8451,g4057);
  IV  NOT_6846(g22198,g19147);
  IV  NOT_6847(g22529,g19549);
  IV  NOT_6848(g34122,I32059);
  IV  NOT_6849(g15799,g13110);
  IV  NOT_6850(I21831,g19127);
  IV  NOT_6851(g13506,g10808);
  IV  NOT_6852(g12088,g7701);
  IV  NOT_6853(g13028,I15650);
  IV  NOT_6854(g20446,g15224);
  IV  NOT_6855(g10386,g6982);
  IV  NOT_6856(g29194,I27492);
  IV  NOT_6857(g9915,g2583);
  IV  NOT_6858(g12860,g10368);
  IV  NOT_6859(g22528,g19801);
  IV  NOT_6860(g6850,g2704);
  IV  NOT_6861(g14386,I16544);
  IV  NOT_6862(g23769,g19074);
  IV  NOT_6863(I11980,g66);
  IV  NOT_6864(g22330,g19801);
  IV  NOT_6865(I13889,g7598);
  IV  NOT_6866(g25542,g22763);
  IV  NOT_6867(g7802,g324);
  IV  NOT_6868(g20059,g17302);
  IV  NOT_6869(g32613,g30673);
  IV  NOT_6870(g8146,g1760);
  IV  NOT_6871(g10096,g5767);
  IV  NOT_6872(g20025,g17271);
  IV  NOT_6873(g8346,g3845);
  IV  NOT_6874(g24059,g21193);
  IV  NOT_6875(g33454,I30980);
  IV  NOT_6876(g14096,I16328);
  IV  NOT_6877(g24025,g21256);
  IV  NOT_6878(g9214,g617);
  IV  NOT_6879(g17529,g15039);
  IV  NOT_6880(g20540,g16646);
  IV  NOT_6881(g12497,g9780);
  IV  NOT_6882(g30292,g28736);
  IV  NOT_6883(I16898,g10615);
  IV  NOT_6884(g23768,g18997);
  IV  NOT_6885(I12884,g4213);
  IV  NOT_6886(I22467,g19662);
  IV  NOT_6887(g20058,g16782);
  IV  NOT_6888(g24540,g22942);
  IV  NOT_6889(g33712,I31561);
  IV  NOT_6890(I26356,g26843);
  IV  NOT_6891(I18307,g12977);
  IV  NOT_6892(g32947,g31376);
  IV  NOT_6893(g19531,g16816);
  IV  NOT_6894(g24058,g20982);
  IV  NOT_6895(g22869,g20875);
  IV  NOT_6896(g17528,g14940);
  IV  NOT_6897(g7558,I12041);
  IV  NOT_6898(g32605,g30614);
  IV  NOT_6899(g8696,g3347);
  IV  NOT_6900(g34409,g34145);
  IV  NOT_6901(I21722,g19264);
  IV  NOT_6902(g22868,g20453);
  IV  NOT_6903(I16521,g10430);
  IV  NOT_6904(g17764,I18758);
  IV  NOT_6905(I12666,g4040);
  IV  NOT_6906(g10429,g7148);
  IV  NOT_6907(g11927,g10207);
  IV  NOT_6908(g23881,g19277);
  IV  NOT_6909(g10857,g8712);
  IV  NOT_6910(g32812,g30825);
  IV  NOT_6911(g25073,I24237);
  IV  NOT_6912(g32463,g31566);
  IV  NOT_6913(g16100,I17471);
  IV  NOT_6914(I32446,g34127);
  IV  NOT_6915(g19676,g17062);
  IV  NOT_6916(g19685,g16987);
  IV  NOT_6917(g31239,g29916);
  IV  NOT_6918(g25274,g22763);
  IV  NOT_6919(g24044,g21127);
  IV  NOT_6920(g16771,g14018);
  IV  NOT_6921(g34408,g34144);
  IV  NOT_6922(I22419,g19638);
  IV  NOT_6923(g19373,g16449);
  IV  NOT_6924(g26575,g25268);
  IV  NOT_6925(g10428,g9631);
  IV  NOT_6926(g32951,g31021);
  IV  NOT_6927(g32972,g31710);
  IV  NOT_6928(g16235,g13437);
  IV  NOT_6929(g32033,g30929);
  IV  NOT_6930(I32059,g33648);
  IV  NOT_6931(g8508,g3827);
  IV  NOT_6932(g19654,g16931);
  IV  NOT_6933(I31361,g33120);
  IV  NOT_6934(g9402,g6209);
  IV  NOT_6935(g9824,g1825);
  IV  NOT_6936(g8944,g370);
  IV  NOT_6937(g8240,g1333);
  IV  NOT_6938(g18661,I19487);
  IV  NOT_6939(g20902,I20870);
  IV  NOT_6940(g18895,g16000);
  IV  NOT_6941(g19800,g17096);
  IV  NOT_6942(I18341,g14308);
  IV  NOT_6943(g19417,g17178);
  IV  NOT_6944(g21662,g16540);
  IV  NOT_6945(g24377,g22594);
  IV  NOT_6946(g7092,g6483);
  IV  NOT_6947(I31500,g33176);
  IV  NOT_6948(g24120,g19984);
  IV  NOT_6949(g23027,g20391);
  IV  NOT_6950(g32795,g31327);
  IV  NOT_6951(g25034,g23695);
  IV  NOT_6952(I23342,g23299);
  IV  NOT_6953(g17709,g14761);
  IV  NOT_6954(g33382,g32033);
  IV  NOT_6955(I12580,g1239);
  IV  NOT_6956(g8443,g3736);
  IV  NOT_6957(g19334,I19818);
  IV  NOT_6958(g20146,g17533);
  IV  NOT_6959(g20738,g15483);
  IV  NOT_6960(I18180,g13605);
  IV  NOT_6961(g25641,I24784);
  IV  NOT_6962(g20562,g17955);
  IV  NOT_6963(g9590,g1882);
  IV  NOT_6964(g21249,g15509);
  IV  NOT_6965(I15981,g11290);
  IV  NOT_6966(g24146,g19422);
  IV  NOT_6967(g6986,g4743);
  IV  NOT_6968(g23249,g21070);
  IV  NOT_6969(I14687,g7753);
  IV  NOT_6970(g11770,I14619);
  IV  NOT_6971(I21199,g17501);
  IV  NOT_6972(I30998,g32453);
  IV  NOT_6973(g20699,g17873);
  IV  NOT_6974(g16515,g13486);
  IV  NOT_6975(g10504,g8763);
  IV  NOT_6976(g11981,I14823);
  IV  NOT_6977(g9657,g2763);
  IV  NOT_6978(g12968,g11793);
  IV  NOT_6979(g17471,g14454);
  IV  NOT_6980(g25153,g23733);
  IV  NOT_6981(I26448,g26860);
  IV  NOT_6982(g8316,g2351);
  IV  NOT_6983(g17087,g14321);
  IV  NOT_6984(g23482,g18833);
  IV  NOT_6985(I25552,g25240);
  IV  NOT_6986(g32514,g30735);
  IV  NOT_6987(I18734,g6373);
  IV  NOT_6988(g24699,g23047);
  IV  NOT_6989(g21248,g15224);
  IV  NOT_6990(g14504,g12361);
  IV  NOT_6991(g19762,g16326);
  IV  NOT_6992(g23248,g20924);
  IV  NOT_6993(g19964,g17200);
  IV  NOT_6994(I22589,g21340);
  IV  NOT_6995(g20698,g17873);
  IV  NOT_6996(g27527,I26195);
  IV  NOT_6997(g25409,g22228);
  IV  NOT_6998(g34575,I32651);
  IV  NOT_6999(I25779,g26424);
  IV  NOT_7000(g32507,g30735);
  IV  NOT_7001(g9556,g5448);
  IV  NOT_7002(I18839,g13716);
  IV  NOT_7003(g23003,I22180);
  IV  NOT_7004(g8565,g3802);
  IV  NOT_7005(g21204,g15656);
  IV  NOT_7006(g33637,I31466);
  IV  NOT_7007(g29177,g27937);
  IV  NOT_7008(g30327,I28582);
  IV  NOT_7009(g33935,I31817);
  IV  NOT_7010(g34711,g34559);
  IV  NOT_7011(g12870,g10374);
  IV  NOT_7012(I11860,g43);
  IV  NOT_7013(g25136,g22457);
  IV  NOT_7014(g34327,g34108);
  IV  NOT_7015(I18667,g6661);
  IV  NOT_7016(I18694,g5666);
  IV  NOT_7017(g32421,g31213);
  IV  NOT_7018(I23330,g22658);
  IV  NOT_7019(I23393,g23414);
  IV  NOT_7020(g10129,g5352);
  IV  NOT_7021(I29441,g30917);
  IV  NOT_7022(g11845,I14663);
  IV  NOT_7023(g9064,g4983);
  IV  NOT_7024(I18131,g13350);
  IV  NOT_7025(g8681,g763);
  IV  NOT_7026(g10002,g6195);
  IV  NOT_7027(I25786,g26424);
  IV  NOT_7028(g10057,g6455);
  IV  NOT_7029(g9899,g6513);
  IV  NOT_7030(I32645,g34367);
  IV  NOT_7031(g7262,g5723);
  IV  NOT_7032(g24366,g22594);
  IV  NOT_7033(g20632,g15171);
  IV  NOT_7034(I15633,g12074);
  IV  NOT_7035(I32699,g34569);
  IV  NOT_7036(I33273,g34984);
  IV  NOT_7037(g30606,I28866);
  IV  NOT_7038(g8697,g3694);
  IV  NOT_7039(I33106,g34855);
  IV  NOT_7040(I14668,g7753);
  IV  NOT_7041(I25356,g24374);
  IV  NOT_7042(g19543,g16349);
  IV  NOT_7043(g30303,g28786);
  IV  NOT_7044(g8914,g4264);
  IV  NOT_7045(I19796,g17870);
  IV  NOT_7046(g17602,g14962);
  IV  NOT_7047(g12867,g10375);
  IV  NOT_7048(g12894,g10401);
  IV  NOT_7049(I17401,g13394);
  IV  NOT_7050(g16584,g13920);
  IV  NOT_7051(g17774,g14902);
  IV  NOT_7052(g23647,g18833);
  IV  NOT_7053(g18889,g15509);
  IV  NOT_7054(g17955,I18865);
  IV  NOT_7055(g18980,g16136);
  IV  NOT_7056(g32541,g30673);
  IV  NOT_7057(g7623,I12103);
  IV  NOT_7058(g10323,I13744);
  IV  NOT_7059(g23945,g21611);
  IV  NOT_7060(g16206,g13437);
  IV  NOT_7061(I25380,g24481);
  IV  NOT_7062(g18095,I18891);
  IV  NOT_7063(g23356,g21070);
  IV  NOT_7064(g32473,g31070);
  IV  NOT_7065(I31463,g33318);
  IV  NOT_7066(g19908,g16540);
  IV  NOT_7067(g22171,g18882);
  IV  NOT_7068(g13191,I15788);
  IV  NOT_7069(g26840,I25562);
  IV  NOT_7070(g20661,g15171);
  IV  NOT_7071(I12654,g1585);
  IV  NOT_7072(g21380,g17955);
  IV  NOT_7073(g10533,g8795);
  IV  NOT_7074(g20547,g15224);
  IV  NOT_7075(g23999,g21468);
  IV  NOT_7076(g32789,g30735);
  IV  NOT_7077(g18888,g15426);
  IV  NOT_7078(g23380,g20619);
  IV  NOT_7079(g33729,I31586);
  IV  NOT_7080(I18443,g13027);
  IV  NOT_7081(g19569,g16349);
  IV  NOT_7082(I14424,g4005);
  IV  NOT_7083(I14016,g9104);
  IV  NOT_7084(I17118,g14363);
  IV  NOT_7085(g16725,g13963);
  IV  NOT_7086(I22748,g19458);
  IV  NOT_7087(g13521,g11357);
  IV  NOT_7088(g22994,g20436);
  IV  NOT_7089(g34982,I33246);
  IV  NOT_7090(g32788,g31327);
  IV  NOT_7091(g32724,g30735);
  IV  NOT_7092(g19747,g17015);
  IV  NOT_7093(g23233,g21037);
  IV  NOT_7094(g21182,g15509);
  IV  NOT_7095(g6789,I11635);
  IV  NOT_7096(g11832,g8011);
  IV  NOT_7097(g23182,g21389);
  IV  NOT_7098(g20715,g15277);
  IV  NOT_7099(g23651,g20655);
  IV  NOT_7100(g32829,g30937);
  IV  NOT_7101(g28080,I26581);
  IV  NOT_7102(g32920,g30825);
  IV  NOT_7103(I18469,g13809);
  IV  NOT_7104(g32535,g31554);
  IV  NOT_7105(g25327,g22161);
  IV  NOT_7106(g32434,g31189);
  IV  NOT_7107(I14830,g10141);
  IV  NOT_7108(I21258,g16540);
  IV  NOT_7109(g24481,I23684);
  IV  NOT_7110(I14893,g9819);
  IV  NOT_7111(g25109,g23666);
  IV  NOT_7112(g12818,g8792);
  IV  NOT_7113(g20551,g17302);
  IV  NOT_7114(g20572,g15833);
  IV  NOT_7115(g9194,g827);
  IV  NOT_7116(g32828,g31710);
  IV  NOT_7117(g18931,g16031);
  IV  NOT_7118(g6987,g4754);
  IV  NOT_7119(g32946,g31327);
  IV  NOT_7120(g10232,g4527);
  IV  NOT_7121(I17276,g13605);
  IV  NOT_7122(g7285,g4643);
  IV  NOT_7123(g11861,g8070);
  IV  NOT_7124(g22919,g21163);
  IV  NOT_7125(g16744,I17964);
  IV  NOT_7126(I17704,g13144);
  IV  NOT_7127(g12978,I15593);
  IV  NOT_7128(g14232,g11083);
  IV  NOT_7129(g9731,g5366);
  IV  NOT_7130(g23331,g20905);
  IV  NOT_7131(I13968,g7697);
  IV  NOT_7132(I32547,g34397);
  IV  NOT_7133(g19751,g16044);
  IV  NOT_7134(I24839,g24298);
  IV  NOT_7135(g9489,g2303);
  IV  NOT_7136(g19772,g17183);
  IV  NOT_7137(g25283,g22763);
  IV  NOT_7138(g34840,I33056);
  IV  NOT_7139(g20127,I20388);
  IV  NOT_7140(I22177,g21366);
  IV  NOT_7141(g23449,g18833);
  IV  NOT_7142(g26483,I25359);
  IV  NOT_7143(g28753,I27235);
  IV  NOT_7144(g9557,g5499);
  IV  NOT_7145(g13926,I16217);
  IV  NOT_7146(g24127,g19984);
  IV  NOT_7147(g13045,g11941);
  IV  NOT_7148(g10261,g4555);
  IV  NOT_7149(I17808,g13311);
  IV  NOT_7150(g9071,g2831);
  IV  NOT_7151(g26862,I25598);
  IV  NOT_7152(g11388,I14395);
  IV  NOT_7153(g23897,g19210);
  IV  NOT_7154(g13099,I15732);
  IV  NOT_7155(g11324,g7542);
  IV  NOT_7156(g23448,g21611);
  IV  NOT_7157(g23961,g19074);
  IV  NOT_7158(g32682,g30825);
  IV  NOT_7159(g24490,g22594);
  IV  NOT_7160(I14705,g7717);
  IV  NOT_7161(g19638,g17324);
  IV  NOT_7162(I17101,g14338);
  IV  NOT_7163(g34192,g33921);
  IV  NOT_7164(I21810,g20596);
  IV  NOT_7165(I16629,g11987);
  IV  NOT_7166(g16652,g13892);
  IV  NOT_7167(g17010,I18138);
  IV  NOT_7168(g23505,g21514);
  IV  NOT_7169(I27543,g28187);
  IV  NOT_7170(g26326,g24872);
  IV  NOT_7171(g8922,I12907);
  IV  NOT_7172(g20385,g18008);
  IV  NOT_7173(I14679,g9332);
  IV  NOT_7174(g13251,I15814);
  IV  NOT_7175(I23375,g23403);
  IV  NOT_7176(g13272,I15837);
  IV  NOT_7177(g19416,g15885);
  IV  NOT_7178(g20103,g17433);
  IV  NOT_7179(g7424,g2465);
  IV  NOT_7180(g24376,g22722);
  IV  NOT_7181(g24385,g22908);
  IV  NOT_7182(g34522,g34271);
  IV  NOT_7183(g7809,g4864);
  IV  NOT_7184(I18143,g13350);
  IV  NOT_7185(g24103,g21209);
  IV  NOT_7186(g23026,g20391);
  IV  NOT_7187(g18088,g13267);
  IV  NOT_7188(g24980,g22384);
  IV  NOT_7189(I16246,g3983);
  IV  NOT_7190(I30971,g32015);
  IV  NOT_7191(I12117,g586);
  IV  NOT_7192(g24095,g21209);
  IV  NOT_7193(g26702,g25309);
  IV  NOT_7194(g17599,g14794);
  IV  NOT_7195(I12000,g582);
  IV  NOT_7196(g25174,g23890);
  IV  NOT_7197(g28696,g27858);
  IV  NOT_7198(g31653,g29713);
  IV  NOT_7199(g6991,g4888);
  IV  NOT_7200(g33653,I31486);
  IV  NOT_7201(I14939,g10216);
  IV  NOT_7202(g7231,g5);
  IV  NOT_7203(g20671,g15509);
  IV  NOT_7204(I17733,g14844);
  IV  NOT_7205(g27018,I25750);
  IV  NOT_7206(g31138,g29778);
  IV  NOT_7207(g32760,g30735);
  IV  NOT_7208(g17086,g14297);
  IV  NOT_7209(g24181,I23387);
  IV  NOT_7210(g7523,g305);
  IV  NOT_7211(g19579,g16000);
  IV  NOT_7212(g22159,I21744);
  IV  NOT_7213(g29941,g28900);
  IV  NOT_7214(g13140,g10632);
  IV  NOT_7215(g7643,g4322);
  IV  NOT_7216(I21792,g21308);
  IV  NOT_7217(I12568,g5005);
  IV  NOT_7218(g12018,g9538);
  IV  NOT_7219(I22009,g21269);
  IV  NOT_7220(g34553,I32621);
  IV  NOT_7221(g10499,I13872);
  IV  NOT_7222(I22665,g21308);
  IV  NOT_7223(I13581,g6727);
  IV  NOT_7224(I18168,g13191);
  IV  NOT_7225(I24278,g23440);
  IV  NOT_7226(I14267,g7835);
  IV  NOT_7227(g32506,g31376);
  IV  NOT_7228(g8784,I12764);
  IV  NOT_7229(I31724,g33076);
  IV  NOT_7230(g33636,I31463);
  IV  NOT_7231(g29185,I27481);
  IV  NOT_7232(I32956,g34654);
  IV  NOT_7233(g30326,I28579);
  IV  NOT_7234(g21723,I21288);
  IV  NOT_7235(g29092,g27800);
  IV  NOT_7236(I32297,g34059);
  IV  NOT_7237(g34949,g34939);
  IV  NOT_7238(g10498,g7161);
  IV  NOT_7239(I32103,g33661);
  IV  NOT_7240(g34326,g34091);
  IV  NOT_7241(g13061,g10981);
  IV  NOT_7242(I31829,g33454);
  IV  NOT_7243(I18479,g13041);
  IV  NOT_7244(g31852,g29385);
  IV  NOT_7245(g6959,g4420);
  IV  NOT_7246(I31535,g33377);
  IV  NOT_7247(g30040,g29025);
  IV  NOT_7248(I13202,g5105);
  IV  NOT_7249(g19586,g16349);
  IV  NOT_7250(I12123,g758);
  IV  NOT_7251(g17125,I18177);
  IV  NOT_7252(g17532,I18479);
  IV  NOT_7253(g27402,I26100);
  IV  NOT_7254(g34536,I32601);
  IV  NOT_7255(I17166,g14536);
  IV  NOT_7256(g28161,I26676);
  IV  NOT_7257(g7634,I12123);
  IV  NOT_7258(g15758,I17276);
  IV  NOT_7259(g21387,I21115);
  IV  NOT_7260(I22485,g21308);
  IV  NOT_7261(I29221,g30307);
  IV  NOT_7262(g23433,g21562);
  IV  NOT_7263(I28419,g29195);
  IV  NOT_7264(I13979,g7733);
  IV  NOT_7265(I32824,g34475);
  IV  NOT_7266(g24426,g22722);
  IV  NOT_7267(g8479,g3057);
  IV  NOT_7268(g20190,g16971);
  IV  NOT_7269(g22144,g18997);
  IV  NOT_7270(I24038,g22202);
  IV  NOT_7271(g23620,I22769);
  IV  NOT_7272(g28709,I27192);
  IV  NOT_7273(g10080,g1982);
  IV  NOT_7274(I17008,g12857);
  IV  NOT_7275(I32671,g34388);
  IV  NOT_7276(g8840,g4277);
  IV  NOT_7277(g9212,g6466);
  IV  NOT_7278(g12866,g10369);
  IV  NOT_7279(I21918,g21290);
  IV  NOT_7280(I17892,g3325);
  IV  NOT_7281(g21343,g16428);
  IV  NOT_7282(I26925,g27015);
  IV  NOT_7283(g8390,g3385);
  IV  NOT_7284(g32927,g30825);
  IV  NOT_7285(g15345,I17108);
  IV  NOT_7286(g14432,g12311);
  IV  NOT_7287(g17680,g14889);
  IV  NOT_7288(g17144,g14085);
  IV  NOT_7289(g26634,g25317);
  IV  NOT_7290(g26851,I25579);
  IV  NOT_7291(g11447,I14450);
  IV  NOT_7292(g7926,g3423);
  IV  NOT_7293(I15162,g10176);
  IV  NOT_7294(g20546,g18008);
  IV  NOT_7295(g20089,g17533);
  IV  NOT_7296(g23971,g20751);
  IV  NOT_7297(I26378,g26850);
  IV  NOT_7298(g19720,I20130);
  IV  NOT_7299(g20211,g16931);
  IV  NOT_7300(I25369,g24891);
  IV  NOT_7301(g24089,g19890);
  IV  NOT_7302(I19851,g16615);
  IV  NOT_7303(g27597,g26745);
  IV  NOT_7304(g21369,g16285);
  IV  NOT_7305(I33291,g34983);
  IV  NOT_7306(g12077,I14939);
  IV  NOT_7307(g32649,g30673);
  IV  NOT_7308(g25553,g22550);
  IV  NOT_7309(g20088,g17533);
  IV  NOT_7310(I27391,g27929);
  IV  NOT_7311(g8356,g54);
  IV  NOT_7312(I20937,g16967);
  IV  NOT_7313(g9229,g5052);
  IV  NOT_7314(I13094,g2724);
  IV  NOT_7315(g14753,g11317);
  IV  NOT_7316(I33173,g34887);
  IV  NOT_7317(g24088,g21209);
  IV  NOT_7318(g19493,g16349);
  IV  NOT_7319(g24024,g21193);
  IV  NOT_7320(g14342,g12163);
  IV  NOT_7321(g34673,I32803);
  IV  NOT_7322(g34847,I33067);
  IV  NOT_7323(g31609,I29211);
  IV  NOT_7324(g29215,I27561);
  IV  NOT_7325(g10031,I13552);
  IV  NOT_7326(g32648,g30614);
  IV  NOT_7327(g32491,g31566);
  IV  NOT_7328(g32903,g31376);
  IV  NOT_7329(g25326,g22228);
  IV  NOT_7330(g14031,I16289);
  IV  NOT_7331(g9822,g125);
  IV  NOT_7332(g10199,g1968);
  IV  NOT_7333(I11801,g6395);
  IV  NOT_7334(I14455,g10197);
  IV  NOT_7335(g16605,g13955);
  IV  NOT_7336(g11472,g7918);
  IV  NOT_7337(I27579,g28184);
  IV  NOT_7338(I29371,g30325);
  IV  NOT_7339(g12923,I15542);
  IV  NOT_7340(g31608,g29653);
  IV  NOT_7341(g18527,I19345);
  IV  NOT_7342(g20497,g18065);
  IV  NOT_7343(g32604,g31154);
  IV  NOT_7344(g34062,g33711);
  IV  NOT_7345(I28588,g29368);
  IV  NOT_7346(g32755,g31672);
  IV  NOT_7347(I30959,g32021);
  IV  NOT_7348(g10198,I13672);
  IV  NOT_7349(g12300,I15144);
  IV  NOT_7350(g11911,g10022);
  IV  NOT_7351(g16812,g13555);
  IV  NOT_7352(g21412,g15758);
  IV  NOT_7353(g32770,g31710);
  IV  NOT_7354(g34933,g34916);
  IV  NOT_7355(g14198,g12180);
  IV  NOT_7356(g32563,g31554);
  IV  NOT_7357(I32089,g33665);
  IV  NOT_7358(I33134,g34906);
  IV  NOT_7359(g13246,g10939);
  IV  NOT_7360(g20700,g17873);
  IV  NOT_7361(g20659,g17873);
  IV  NOT_7362(g34851,I33075);
  IV  NOT_7363(g20625,g15348);
  IV  NOT_7364(g10393,g6991);
  IV  NOT_7365(g24126,g19935);
  IV  NOT_7366(g24625,g23135);
  IV  NOT_7367(g14330,I16486);
  IV  NOT_7368(g24987,g23630);
  IV  NOT_7369(g8954,g1079);
  IV  NOT_7370(g7543,I12033);
  IV  NOT_7371(g31799,g29385);
  IV  NOT_7372(g23896,g19210);
  IV  NOT_7373(g25564,g22312);
  IV  NOT_7374(g8363,g239);
  IV  NOT_7375(g18894,g16000);
  IV  NOT_7376(g31813,g29385);
  IV  NOT_7377(g21228,g17531);
  IV  NOT_7378(g33799,g33299);
  IV  NOT_7379(g10365,g6867);
  IV  NOT_7380(g22224,g19277);
  IV  NOT_7381(g33813,I31659);
  IV  NOT_7382(g8032,I12355);
  IV  NOT_7383(g19517,g16777);
  IV  NOT_7384(g23228,g21070);
  IV  NOT_7385(I18373,g13011);
  IV  NOT_7386(g29906,g28793);
  IV  NOT_7387(g29348,g28194);
  IV  NOT_7388(g16795,I18009);
  IV  NOT_7389(g10960,g9007);
  IV  NOT_7390(I17675,g13394);
  IV  NOT_7391(g23011,g20330);
  IV  NOT_7392(g31798,g29385);
  IV  NOT_7393(g32767,g30735);
  IV  NOT_7394(g32794,g30937);
  IV  NOT_7395(I14623,g8925);
  IV  NOT_7396(g11147,g8417);
  IV  NOT_7397(g11754,g8229);
  IV  NOT_7398(I17154,g13605);
  IV  NOT_7399(I23680,g23219);
  IV  NOT_7400(g25183,g22763);
  IV  NOT_7401(g32899,g31021);
  IV  NOT_7402(g7534,g1367);
  IV  NOT_7403(g31805,g29385);
  IV  NOT_7404(g17224,I18248);
  IV  NOT_7405(g16514,g14139);
  IV  NOT_7406(g12885,g10382);
  IV  NOT_7407(g22495,g19801);
  IV  NOT_7408(g17308,g14876);
  IV  NOT_7409(g23582,I22729);
  IV  NOT_7410(g32633,g31154);
  IV  NOT_7411(g32898,g30825);
  IV  NOT_7412(I32659,g34391);
  IV  NOT_7413(g15048,I16969);
  IV  NOT_7414(g9620,g6187);
  IV  NOT_7415(g9462,g6215);
  IV  NOT_7416(I23336,g22721);
  IV  NOT_7417(I19756,g17812);
  IV  NOT_7418(g19362,g16072);
  IV  NOT_7419(g7927,g4064);
  IV  NOT_7420(g34574,I32648);
  IV  NOT_7421(g32719,g31672);
  IV  NOT_7422(I12041,g2741);
  IV  NOT_7423(g20060,g16540);
  IV  NOT_7424(g34047,g33637);
  IV  NOT_7425(g18979,g16136);
  IV  NOT_7426(g19523,g16100);
  IV  NOT_7427(g24060,g21256);
  IV  NOT_7428(g8912,g4180);
  IV  NOT_7429(I16120,g11868);
  IV  NOT_7430(g33934,I31814);
  IV  NOT_7431(g10708,g7836);
  IV  NOT_7432(g20197,g16987);
  IV  NOT_7433(g6928,I11716);
  IV  NOT_7434(I12746,g4087);
  IV  NOT_7435(g21379,g17873);
  IV  NOT_7436(g34311,g34097);
  IV  NOT_7437(I12493,g5002);
  IV  NOT_7438(g22976,I22149);
  IV  NOT_7439(g22985,g20330);
  IV  NOT_7440(g32718,g30825);
  IV  NOT_7441(g32521,g31376);
  IV  NOT_7442(g10087,I13597);
  IV  NOT_7443(g23925,g21514);
  IV  NOT_7444(g8357,I12538);
  IV  NOT_7445(g18978,g16000);
  IV  NOT_7446(g7946,I12314);
  IV  NOT_7447(g7660,I12144);
  IV  NOT_7448(g29653,I27927);
  IV  NOT_7449(I22729,g21308);
  IV  NOT_7450(g26820,I25534);
  IV  NOT_7451(g21050,g17873);
  IV  NOT_7452(g20527,g18008);
  IV  NOT_7453(I13597,g4417);
  IV  NOT_7454(g11367,I14381);
  IV  NOT_7455(g28918,g27832);
  IV  NOT_7456(g32832,g30735);
  IV  NOT_7457(I20321,g16920);
  IV  NOT_7458(g23378,g21070);
  IV  NOT_7459(g13394,I15915);
  IV  NOT_7460(I31491,g33283);
  IV  NOT_7461(g33761,I31616);
  IV  NOT_7462(g24527,g22670);
  IV  NOT_7463(g7903,g969);
  IV  NOT_7464(g30072,I28301);
  IV  NOT_7465(g17687,g15042);
  IV  NOT_7466(I31604,g33176);
  IV  NOT_7467(g28079,I26578);
  IV  NOT_7468(g10043,g1632);
  IV  NOT_7469(I13280,g6140);
  IV  NOT_7470(g7513,g6315);
  IV  NOT_7471(g26731,g25470);
  IV  NOT_7472(g34592,I32684);
  IV  NOT_7473(I11688,g70);
  IV  NOT_7474(I16698,g12077);
  IV  NOT_7475(g29333,g28167);
  IV  NOT_7476(g16473,g13977);
  IV  NOT_7477(I31770,g33197);
  IV  NOT_7478(g32861,g31376);
  IV  NOT_7479(g9842,g3274);
  IV  NOT_7480(g23944,g19147);
  IV  NOT_7481(g32573,g30825);
  IV  NOT_7482(g18094,I18888);
  IV  NOT_7483(g31013,g29679);
  IV  NOT_7484(I14589,g8818);
  IV  NOT_7485(g25213,g23293);
  IV  NOT_7486(g19437,g16349);
  IV  NOT_7487(g20503,g15373);
  IV  NOT_7488(g9298,g5080);
  IV  NOT_7489(g28598,g27717);
  IV  NOT_7490(I18909,g16873);
  IV  NOT_7491(g9392,g5869);
  IV  NOT_7492(g32926,g31376);
  IV  NOT_7493(I32855,g34540);
  IV  NOT_7494(g7178,g4392);
  IV  NOT_7495(g7436,g5276);
  IV  NOT_7496(I14836,g9688);
  IV  NOT_7497(g8626,g4040);
  IV  NOT_7498(g21681,I21242);
  IV  NOT_7499(g29963,g28931);
  IV  NOT_7500(g16724,g14079);
  IV  NOT_7501(g22842,g19875);
  IV  NOT_7502(g23681,g21012);
  IV  NOT_7503(I18117,g13302);
  IV  NOT_7504(g32612,g30614);
  IV  NOT_7505(g16325,g13223);
  IV  NOT_7506(g18877,g15224);
  IV  NOT_7507(I23309,g21677);
  IV  NOT_7508(g25452,g22228);
  IV  NOT_7509(g15371,I17114);
  IV  NOT_7510(g25047,g23733);
  IV  NOT_7511(g32099,g31009);
  IV  NOT_7512(g10375,g6941);
  IV  NOT_7513(I21288,g18216);
  IV  NOT_7514(g34820,I33034);
  IV  NOT_7515(g16920,I18086);
  IV  NOT_7516(g20714,g15277);
  IV  NOT_7517(g20450,g15277);
  IV  NOT_7518(g23429,g20453);
  IV  NOT_7519(g32701,g31376);
  IV  NOT_7520(g12076,g9280);
  IV  NOT_7521(g7335,g2287);
  IV  NOT_7522(g7831,I12227);
  IV  NOT_7523(I14119,g7824);
  IV  NOT_7524(g32777,g31710);
  IV  NOT_7525(g32534,g30673);
  IV  NOT_7526(g12721,g10061);
  IV  NOT_7527(g34152,I32109);
  IV  NOT_7528(g20707,g18008);
  IV  NOT_7529(g21428,g15758);
  IV  NOT_7530(I22622,g21209);
  IV  NOT_7531(g20910,g15171);
  IV  NOT_7532(g34846,I33064);
  IV  NOT_7533(g23793,g19074);
  IV  NOT_7534(g12054,g7690);
  IV  NOT_7535(g17392,g14924);
  IV  NOT_7536(g19600,g16164);
  IV  NOT_7537(g10337,g5016);
  IV  NOT_7538(g24819,I23998);
  IV  NOT_7539(g19781,g16489);
  IV  NOT_7540(g17489,g12955);
  IV  NOT_7541(I24334,g22976);
  IV  NOT_7542(g20496,g17929);
  IV  NOT_7543(g7805,g4366);
  IV  NOT_7544(g7916,I12300);
  IV  NOT_7545(g25051,I24215);
  IV  NOT_7546(g25072,g23630);
  IV  NOT_7547(g24818,g23191);
  IV  NOT_7548(g32462,g30673);
  IV  NOT_7549(I14749,g10031);
  IV  NOT_7550(g24979,g22369);
  IV  NOT_7551(g21690,g16540);
  IV  NOT_7552(g22830,g20283);
  IV  NOT_7553(g19952,g15915);
  IV  NOT_7554(g24055,g19968);
  IV  NOT_7555(g7749,g996);
  IV  NOT_7556(g19351,g17367);
  IV  NOT_7557(I12523,g3794);
  IV  NOT_7558(g23549,g18833);
  IV  NOT_7559(g27773,I26378);
  IV  NOT_7560(g20070,g16173);
  IV  NOT_7561(g20978,g15595);
  IV  NOT_7562(g24111,g19890);
  IV  NOT_7563(g28656,g27742);
  IV  NOT_7564(g9708,g2741);
  IV  NOT_7565(g24070,g20014);
  IV  NOT_7566(g24978,g22342);
  IV  NOT_7567(g34691,I32843);
  IV  NOT_7568(g29312,g28877);
  IV  NOT_7569(g20590,g15426);
  IV  NOT_7570(g22544,g19589);
  IV  NOT_7571(g22865,g20330);
  IV  NOT_7572(g23548,g18833);
  IV  NOT_7573(g8778,I12758);
  IV  NOT_7574(g29115,g27779);
  IV  NOT_7575(g7947,g1500);
  IV  NOT_7576(I20216,g15862);
  IV  NOT_7577(g24986,g23590);
  IV  NOT_7578(I14305,g8805);
  IV  NOT_7579(g9252,g4304);
  IV  NOT_7580(I26880,g27527);
  IV  NOT_7581(g23504,g21468);
  IV  NOT_7582(g13902,g11389);
  IV  NOT_7583(g13301,g10862);
  IV  NOT_7584(g31771,I29337);
  IV  NOT_7585(g19264,I19802);
  IV  NOT_7586(g18917,g16077);
  IV  NOT_7587(g19790,g16971);
  IV  NOT_7588(g20384,g18008);
  IV  NOT_7589(g12180,g9477);
  IV  NOT_7590(g9958,g6148);
  IV  NOT_7591(g29921,g28864);
  IV  NOT_7592(g13120,g10632);
  IV  NOT_7593(I18293,g1079);
  IV  NOT_7594(g24384,g22885);
  IV  NOT_7595(g25820,g25051);
  IV  NOT_7596(I26512,g26817);
  IV  NOT_7597(I17653,g14276);
  IV  NOT_7598(g20067,g17328);
  IV  NOT_7599(g32766,g31376);
  IV  NOT_7600(g6955,I11726);
  IV  NOT_7601(g29745,g28500);
  IV  NOT_7602(g24067,g21256);
  IV  NOT_7603(g24094,g21143);
  IV  NOT_7604(g11562,g7648);
  IV  NOT_7605(g17713,g12947);
  IV  NOT_7606(I18265,g13350);
  IV  NOT_7607(g34929,I33179);
  IV  NOT_7608(g27930,I26451);
  IV  NOT_7609(I12437,g4999);
  IV  NOT_7610(g27993,I26503);
  IV  NOT_7611(g8075,g3742);
  IV  NOT_7612(g32871,g30937);
  IV  NOT_7613(g30020,g29097);
  IV  NOT_7614(g30928,I28908);
  IV  NOT_7615(g22189,I21769);
  IV  NOT_7616(g8475,I12608);
  IV  NOT_7617(g26105,I25146);
  IV  NOT_7618(g9829,g2250);
  IV  NOT_7619(g12839,g10350);
  IV  NOT_7620(g6814,g632);
  IV  NOT_7621(g12930,g12347);
  IV  NOT_7622(g7873,g1266);
  IV  NOT_7623(g26743,g25476);
  IV  NOT_7624(g26827,g24819);
  IV  NOT_7625(g34583,I32665);
  IV  NOT_7626(g7632,I12117);
  IV  NOT_7627(g34928,I33176);
  IV  NOT_7628(g7095,g6545);
  IV  NOT_7629(I17636,g14252);
  IV  NOT_7630(g21057,g15426);
  IV  NOT_7631(g23002,I22177);
  IV  NOT_7632(g10079,g1950);
  IV  NOT_7633(g11290,I14326);
  IV  NOT_7634(g24150,g19268);
  IV  NOT_7635(g23057,g20453);
  IV  NOT_7636(I28594,g29379);
  IV  NOT_7637(g9911,g2384);
  IV  NOT_7638(g7495,g4375);
  IV  NOT_7639(g14545,g12768);
  IV  NOT_7640(g7437,g5666);
  IV  NOT_7641(g17610,g15008);
  IV  NOT_7642(I27253,g27996);
  IV  NOT_7643(I30995,g32449);
  IV  NOT_7644(g12838,g10353);
  IV  NOT_7645(g23128,g20283);
  IV  NOT_7646(I20569,g16486);
  IV  NOT_7647(I17852,g3625);
  IV  NOT_7648(g10078,g1854);
  IV  NOT_7649(g21245,I20982);
  IV  NOT_7650(g24019,g19968);
  IV  NOT_7651(g17189,g14708);
  IV  NOT_7652(g23245,g20785);
  IV  NOT_7653(I13287,g110);
  IV  NOT_7654(g26769,g25400);
  IV  NOT_7655(g8526,g1526);
  IV  NOT_7656(g19208,g17367);
  IV  NOT_7657(g20695,I20781);
  IV  NOT_7658(I20747,g17141);
  IV  NOT_7659(I31701,g33164);
  IV  NOT_7660(g21299,g16600);
  IV  NOT_7661(g30113,g29154);
  IV  NOT_7662(g9733,g5736);
  IV  NOT_7663(g10086,g2193);
  IV  NOT_7664(g23323,g20283);
  IV  NOT_7665(g23299,I22400);
  IV  NOT_7666(g9974,g2518);
  IV  NOT_7667(I32067,g33661);
  IV  NOT_7668(g17188,I18224);
  IV  NOT_7669(I11721,g4145);
  IV  NOT_7670(g17124,g14051);
  IV  NOT_7671(g17678,I18653);
  IV  NOT_7672(g34787,I32991);
  IV  NOT_7673(g26803,g25389);
  IV  NOT_7674(g12487,g9340);
  IV  NOT_7675(g20526,g15171);
  IV  NOT_7676(I22576,g21282);
  IV  NOT_7677(I28185,g28803);
  IV  NOT_7678(I18835,g6365);
  IV  NOT_7679(I13054,g6744);
  IV  NOT_7680(g24526,g22942);
  IV  NOT_7681(g19542,g16349);
  IV  NOT_7682(g30302,g28924);
  IV  NOT_7683(g7752,g1542);
  IV  NOT_7684(I16181,g3672);
  IV  NOT_7685(g18102,I18912);
  IV  NOT_7686(g8439,g3129);
  IV  NOT_7687(g9073,g150);
  IV  NOT_7688(g32629,g31376);
  IV  NOT_7689(g34302,I32305);
  IV  NOT_7690(I26989,g27277);
  IV  NOT_7691(I32150,g33923);
  IV  NOT_7692(g30105,I28336);
  IV  NOT_7693(g6836,g1322);
  IV  NOT_7694(g7917,g1157);
  IV  NOT_7695(I14630,g7717);
  IV  NOT_7696(g27279,g26330);
  IV  NOT_7697(g32472,g30825);
  IV  NOT_7698(g10159,g4477);
  IV  NOT_7699(g34827,I33041);
  IV  NOT_7700(g10532,g10233);
  IV  NOT_7701(g32628,g31542);
  IV  NOT_7702(g17093,I18165);
  IV  NOT_7703(g6918,g3639);
  IV  NOT_7704(g32911,g31376);
  IV  NOT_7705(g14125,I16345);
  IV  NOT_7706(g15344,g14851);
  IV  NOT_7707(g10158,g2461);
  IV  NOT_7708(g11403,g7595);
  IV  NOT_7709(g11547,I14505);
  IV  NOT_7710(g13895,I16193);
  IV  NOT_7711(g20917,g15224);
  IV  NOT_7712(I33140,g34884);
  IV  NOT_7713(I28883,g30105);
  IV  NOT_7714(g23232,I22331);
  IV  NOT_7715(g24866,I24038);
  IV  NOT_7716(g19905,g15885);
  IV  NOT_7717(I12790,g4340);
  IV  NOT_7718(I17609,g13510);
  IV  NOT_7719(g34769,I32953);
  IV  NOT_7720(I11655,g1246);
  IV  NOT_7721(g18876,g15373);
  IV  NOT_7722(g18885,g15979);
  IV  NOT_7723(g10353,g6803);
  IV  NOT_7724(g25046,g23729);
  IV  NOT_7725(g6993,g4859);
  IV  NOT_7726(g10295,I13723);
  IV  NOT_7727(g8919,I12896);
  IV  NOT_7728(g21697,I21258);
  IV  NOT_7729(g29013,I27368);
  IV  NOT_7730(I29981,g31591);
  IV  NOT_7731(g34768,I32950);
  IV  NOT_7732(g12039,I14899);
  IV  NOT_7733(g13715,g10573);
  IV  NOT_7734(I22745,g19458);
  IV  NOT_7735(g29214,I27558);
  IV  NOT_7736(g27038,g25932);
  IV  NOT_7737(g9206,g5164);
  IV  NOT_7738(g32591,g30614);
  IV  NOT_7739(I15572,g10499);
  IV  NOT_7740(g23995,g19277);
  IV  NOT_7741(g32776,g31672);
  IV  NOT_7742(g32785,g31710);
  IV  NOT_7743(I30989,g32441);
  IV  NOT_7744(g19565,g16000);
  IV  NOT_7745(g24077,g20720);
  IV  NOT_7746(g20706,g18008);
  IV  NOT_7747(I11734,g4473);
  IV  NOT_7748(g23880,g19210);
  IV  NOT_7749(g12038,I14896);
  IV  NOT_7750(g20597,g17847);
  IV  NOT_7751(I21042,g15824);
  IV  NOT_7752(g32754,g30825);
  IV  NOT_7753(I14570,g7932);
  IV  NOT_7754(g33435,I30959);
  IV  NOT_7755(g25282,g22763);
  IV  NOT_7756(I21189,g17475);
  IV  NOT_7757(g14336,I16498);
  IV  NOT_7758(g27187,I25882);
  IV  NOT_7759(g7296,g5313);
  IV  NOT_7760(g23512,g20248);
  IV  NOT_7761(g8616,g2803);
  IV  NOT_7762(g28752,I27232);
  IV  NOT_7763(g20923,g15277);
  IV  NOT_7764(g27975,g26694);
  IV  NOT_7765(g32859,g30614);
  IV  NOT_7766(g32825,g30735);
  IV  NOT_7767(g32950,g31672);
  IV  NOT_7768(g28954,g27830);
  IV  NOT_7769(g26710,g25349);
  IV  NOT_7770(g18660,I19484);
  IV  NOT_7771(g20624,g18065);
  IV  NOT_7772(g22455,g19801);
  IV  NOT_7773(g12975,g12752);
  IV  NOT_7774(g7532,g1157);
  IV  NOT_7775(I13694,g117);
  IV  NOT_7776(I16024,g11171);
  IV  NOT_7777(g32858,g31327);
  IV  NOT_7778(g33744,I31604);
  IV  NOT_7779(g7553,g1274);
  IV  NOT_7780(g8404,g5005);
  IV  NOT_7781(g15506,I17131);
  IV  NOT_7782(g31849,g29385);
  IV  NOT_7783(g8647,g3416);
  IV  NOT_7784(g14631,g12239);
  IV  NOT_7785(g10364,g6869);
  IV  NOT_7786(g19409,g16431);
  IV  NOT_7787(I14567,g9708);
  IV  NOT_7788(g12143,I14999);
  IV  NOT_7789(g20102,g17533);
  IV  NOT_7790(g16767,I17989);
  IV  NOT_7791(g20157,g16886);
  IV  NOT_7792(g25640,I24781);
  IV  NOT_7793(g12937,g12419);
  IV  NOT_7794(g28669,g27705);
  IV  NOT_7795(g26081,g24619);
  IV  NOT_7796(g8764,g4826);
  IV  NOT_7797(g22201,g19277);
  IV  NOT_7798(g24102,g21143);
  IV  NOT_7799(g23445,I22564);
  IV  NOT_7800(g31848,g29385);
  IV  NOT_7801(g18916,g16053);
  IV  NOT_7802(g24157,I23315);
  IV  NOT_7803(g32844,g30937);
  IV  NOT_7804(g9898,g6444);
  AN2 AND2_0(g33848,g33261,g20384);
  AN2 AND2_1(g28260,g27703,g26518);
  AN2 AND2_2(g17617,g7885,g13326);
  AN2 AND2_3(g18550,g2819,g15277);
  AN2 AND2_4(g25768,g2912,g24560);
  AN2 AND2_5(g25803,g24798,g21024);
  AN2 AND2_6(g31141,g12224,g30038);
  AN3 AND3_0(I26960,g24995,g26424,g22698);
  AN2 AND2_7(g22075,g6247,g19210);
  AN2 AND2_8(g18314,g1585,g16931);
  AN2 AND2_9(g33652,g33393,g18889);
  AN2 AND2_10(g18287,g1442,g16449);
  AN2 AND2_11(g27410,g26549,g17527);
  AN2 AND2_12(g16633,g5196,g14921);
  AN2 AND2_13(g30248,g28743,g23938);
  AN2 AND2_14(g34482,g34405,g18917);
  AN2 AND2_15(g23498,g20234,g12998);
  AN2 AND2_16(g28489,g27010,g12417);
  AN2 AND2_17(g26356,g15581,g25523);
  AN2 AND2_18(g18307,g1559,g16931);
  AN2 AND2_19(g29771,g28322,g23242);
  AN2 AND2_20(g30003,g28149,g9021);
  AN2 AND2_21(g34710,g34553,g20903);
  AN2 AND2_22(g16191,g5475,g14262);
  AN2 AND2_23(g22623,g19337,g19470);
  AN2 AND2_24(g21989,g5587,g19074);
  AN2 AND2_25(g30204,g28670,g23868);
  AN2 AND2_26(g13671,g4498,g10532);
  AN2 AND2_27(g26826,g24907,g15747);
  AN2 AND2_28(g27666,g26865,g23521);
  AN4 AND4_0(I31246,g31672,g31839,g32810,g32811);
  AN2 AND2_29(g18721,g15138,g16077);
  AN2 AND2_30(g22037,g5941,g19147);
  AN2 AND2_31(g25881,g3821,g24685);
  AN2 AND2_32(g26380,g19572,g25547);
  AN2 AND2_33(g33263,g32393,g25481);
  AN2 AND2_34(g18596,g2941,g16349);
  AN2 AND2_35(g32420,g31127,g19533);
  AN2 AND2_36(g28488,g27969,g17713);
  AN2 AND2_37(g27363,g10231,g26812);
  AN2 AND2_38(g23056,g16052,g19860);
  AN3 AND3_1(g27217,g26236,g8418,g2610);
  AN2 AND2_39(g29683,g1821,g29046);
  AN2 AND2_40(g18243,g1189,g16431);
  AN2 AND2_41(g33332,g32217,g20608);
  AN3 AND3_2(I17692,g14988,g11450,g6756);
  AN2 AND2_42(g21988,g5583,g19074);
  AN2 AND2_43(g26090,g1624,g25081);
  AN2 AND2_44(g21924,g5057,g21468);
  AN2 AND2_45(g28558,g7301,g27046);
  AN2 AND2_46(g18431,g2185,g18008);
  AN2 AND2_47(g26233,g2279,g25309);
  AN4 AND4_1(I31071,g31170,g31808,g32557,g32558);
  AN2 AND2_48(g26182,g9978,g25317);
  AN2 AND2_49(g26651,g22707,g24425);
  AN2 AND2_50(g12015,g1002,g7567);
  AN2 AND2_51(g34081,g33706,g19552);
  AN2 AND2_52(g27486,g26519,g17645);
  AN2 AND2_53(g31962,g8033,g31013);
  AN2 AND2_54(g24763,g17569,g22457);
  AN2 AND2_55(g33406,g32355,g21399);
  AN2 AND2_56(g18269,g15069,g16031);
  AN2 AND2_57(g33361,g32257,g20911);
  AN2 AND2_58(g15903,g13796,g13223);
  AN2 AND2_59(g18773,g5694,g15615);
  AN4 AND4_2(I31147,g32668,g32669,g32670,g32671);
  AN2 AND2_60(g18341,g1648,g17873);
  AN2 AND2_61(g29515,g28888,g22342);
  AN2 AND2_62(g29882,g2361,g29151);
  AN2 AND2_63(g18268,g1280,g16000);
  AN2 AND2_64(g29991,g29179,g12922);
  AN2 AND2_65(g21753,g3179,g20785);
  AN2 AND2_66(g31500,g29802,g23449);
  AN2 AND2_67(g18156,g572,g17533);
  AN2 AND2_68(g18655,g15106,g14454);
  AN3 AND3_3(g33500,g32744,I31196,I31197);
  AN2 AND2_69(g24660,g22648,g19737);
  AN2 AND2_70(g33833,g33093,g25852);
  AN2 AND2_71(g32203,g4249,g31327);
  AN2 AND2_72(g18180,g767,g17328);
  AN2 AND2_73(g26513,g19501,g24365);
  AN2 AND2_74(g17418,g9618,g14407);
  AN3 AND3_4(I27409,g25556,g26424,g22698);
  AN2 AND2_75(g34999,g34998,g23085);
  AN2 AND2_76(g18670,g4621,g15758);
  AN2 AND2_77(g34380,g34158,g20571);
  AN3 AND3_5(g25482,g5752,g23816,I24597);
  AN2 AND2_78(g32044,g31483,g20085);
  AN4 AND4_3(I24684,g20014,g24033,g24034,g24035);
  AN2 AND2_79(g16612,g5603,g14927);
  AN2 AND2_80(g21736,g3065,g20330);
  AN2 AND2_81(g11546,g7289,g4375);
  AN2 AND2_82(g21887,g15101,g19801);
  AN2 AND2_83(g30233,g28720,g23913);
  AN2 AND2_84(g18734,g4966,g16826);
  AN4 AND4_4(I31151,g30825,g31822,g32673,g32674);
  AN2 AND2_85(g16324,g13657,g182);
  AN4 AND4_5(I31172,g32703,g32704,g32705,g32706);
  AN2 AND2_86(g18335,g1687,g17873);
  AN2 AND2_87(g16701,g5547,g14845);
  AN2 AND2_88(g22589,g19267,g19451);
  AN2 AND2_89(g32281,g31257,g20500);
  AN2 AND2_90(g34182,g33691,g24384);
  AN2 AND2_91(g28255,g8515,g27983);
  AN2 AND2_92(g16534,g5575,g14665);
  AN2 AND2_93(g28679,g27572,g20638);
  AN2 AND2_94(g11024,g5436,g9070);
  AN2 AND2_95(g16098,g5148,g14238);
  AN3 AND3_6(I13937,g7340,g7293,g7261);
  AN2 AND2_96(g18993,g11224,g16172);
  AN2 AND2_97(g24550,g3684,g23308);
  AN2 AND2_98(g32301,g31276,g20547);
  AN2 AND2_99(g14643,g11998,g12023);
  AN2 AND2_100(g24314,g4515,g22228);
  AN2 AND2_101(g22588,g79,g20078);
  AN2 AND2_102(g21843,g3869,g21070);
  AN2 AND2_103(g32120,g31639,g29941);
  AN2 AND2_104(g24287,g4401,g22550);
  AN2 AND2_105(g28124,g27368,g22842);
  AN2 AND2_106(g15794,g3239,g14008);
  AN2 AND2_107(g18667,g4601,g17367);
  AN2 AND2_108(g18694,g4722,g16053);
  AN2 AND2_109(g12179,g9745,g10027);
  AN2 AND2_110(g24307,g4486,g22228);
  AN2 AND2_111(g29584,g1706,g29018);
  AN2 AND2_112(g27178,g25997,g16652);
  AN2 AND2_113(g21764,g3227,g20785);
  AN2 AND2_114(g11497,g6398,g7192);
  AN2 AND2_115(g18131,g482,g16971);
  AN3 AND3_7(g29206,g24124,I27528,I27529);
  AN2 AND2_116(g13497,g2724,g12155);
  AN2 AND2_117(g28686,g27574,g20650);
  AN2 AND2_118(g32146,g31624,g29978);
  AN4 AND4_6(g28939,g17321,g25184,g26424,g27421);
  AN2 AND2_119(g24721,g17488,g22369);
  AN2 AND2_120(g22119,g6581,g19277);
  AN2 AND2_121(g21869,g4087,g19801);
  AN3 AND3_8(g27186,g26195,g8316,g2342);
  AN2 AND2_122(g31273,g30143,g27779);
  AN2 AND2_123(g34513,g9003,g34346);
  AN2 AND2_124(g21960,g5421,g21514);
  AN2 AND2_125(g27676,g26377,g20627);
  AN2 AND2_126(g27685,g13032,g25895);
  AN2 AND2_127(g15633,g3841,g13584);
  AN2 AND2_128(g33106,g32408,g18990);
  AN2 AND2_129(g18487,g2441,g15426);
  AN2 AND2_130(g27373,g26488,g17477);
  AN2 AND2_131(g29759,g28308,g23226);
  AN2 AND2_132(g22118,g6605,g19277);
  AN2 AND2_133(g32290,g31267,g20525);
  AN2 AND2_134(g11126,g6035,g10185);
  AN2 AND2_135(g12186,g1178,g7519);
  AN3 AND3_9(g28267,g7328,g2227,g27421);
  AN2 AND2_136(g17401,g1083,g13143);
  AN2 AND2_137(g21868,g4076,g19801);
  AN2 AND2_138(g18619,g3466,g17062);
  AN2 AND2_139(g18502,g2567,g15509);
  AN2 AND2_140(g22022,g5873,g19147);
  AN2 AND2_141(g34961,g34944,g23019);
  AN2 AND2_142(g12953,g411,g11048);
  AN2 AND2_143(g18557,g2771,g15277);
  AN3 AND3_10(g33812,g23088,g33187,g9104);
  AN2 AND2_144(g18210,g936,g15938);
  AN2 AND2_145(g29758,g28306,g23222);
  AN2 AND2_146(g17119,g5272,g14800);
  AN3 AND3_11(g33463,g32477,I31011,I31012);
  AN4 AND4_7(I31227,g32784,g32785,g32786,g32787);
  AN2 AND2_147(g18618,g3457,g17062);
  AN2 AND2_148(g18443,g2265,g18008);
  AN2 AND2_149(g24773,g22832,g19872);
  AN2 AND2_150(g21709,g283,g20283);
  AN2 AND2_151(g18279,g1361,g16136);
  AN2 AND2_152(g30026,g28476,g25064);
  AN2 AND2_153(g33371,g32280,g21155);
  AN2 AND2_154(g30212,g28687,g23879);
  AN2 AND2_155(g16766,g6649,g12915);
  AN2 AND2_156(g26387,g24813,g20231);
  AN2 AND2_157(g27334,g12539,g26769);
  AN2 AND2_158(g34212,g33761,g22689);
  AN2 AND2_159(g28219,g9316,g27573);
  AN2 AND2_160(g21708,g15049,g20283);
  AN2 AND2_161(g18278,g1345,g16136);
  AN3 AND3_12(I16111,g8691,g11409,g11381);
  AN4 AND4_8(g26148,g25357,g11724,g11709,g11686);
  AN2 AND2_162(g23708,g19050,g9104);
  AN2 AND2_163(g16871,g6597,g14908);
  AN2 AND2_164(g29345,g4749,g28376);
  AN2 AND2_165(g22053,g6116,g21611);
  AN2 AND2_166(g23471,g20148,g20523);
  AN2 AND2_167(g26097,g5821,g25092);
  AN2 AND2_168(g18469,g2399,g15224);
  AN2 AND2_169(g24670,g5138,g23590);
  AN2 AND2_170(g33795,g33138,g20782);
  AN2 AND2_171(g28218,g27768,g26645);
  AN2 AND2_172(g29940,g1740,g28758);
  AN2 AND2_173(g26104,g2250,g25101);
  AN2 AND2_174(g18286,g1404,g16164);
  AN2 AND2_175(g22900,g17137,g19697);
  AN4 AND4_9(g27762,g22472,g25226,g26424,g26218);
  AN2 AND2_176(g15861,g3957,g14170);
  AN2 AND2_177(g8690,g2941,g2936);
  AN2 AND2_178(g27964,g25956,g22492);
  AN2 AND2_179(g18468,g2393,g15224);
  AN3 AND3_13(g25331,g5366,g22194,I24508);
  AN2 AND2_180(g18306,g15074,g16931);
  AN2 AND2_181(g12762,g4358,g8977);
  AN2 AND2_182(g22036,g5937,g19147);
  AN2 AND2_183(g25449,g6946,g22496);
  AN2 AND2_184(g13060,g8587,g11110);
  AN2 AND2_185(g31514,g20041,g29956);
  AN2 AND2_186(g32403,g31117,g15842);
  AN2 AND2_187(g27216,g26055,g16725);
  AN3 AND3_14(g33514,g32844,I31266,I31267);
  AN2 AND2_188(g22101,g6474,g18833);
  AN2 AND2_189(g24930,g4826,g23948);
  AN2 AND2_190(g29652,g2667,g29157);
  AN2 AND2_191(g29804,g1592,g29014);
  AN2 AND2_192(g17809,g7873,g13125);
  AN4 AND4_10(I31281,g30735,g31845,g32861,g32862);
  AN2 AND2_193(g28160,g26309,g27463);
  AN2 AND2_194(g15612,g3143,g13530);
  AN2 AND2_195(g25448,g11202,g22680);
  AN2 AND2_196(g18815,g6523,g15483);
  AN2 AND2_197(g30149,g28605,g21248);
  AN2 AND2_198(g25961,g25199,g20682);
  AN3 AND3_15(I27381,g25549,g26424,g22698);
  AN3 AND3_16(g33507,g32795,I31231,I31232);
  AN4 AND4_11(I31301,g31327,g31849,g32889,g32890);
  AN2 AND2_199(g20131,g15170,g14309);
  AN2 AND2_200(g15701,g3821,g13584);
  AN3 AND3_17(g10705,g6850,g10219,g2689);
  AN2 AND2_201(g18601,g3106,g16987);
  AN2 AND2_202(g13411,g4955,g11834);
  AN2 AND2_203(g18187,g794,g17328);
  AN2 AND2_204(g18677,g4639,g15758);
  AN2 AND2_205(g14610,g1484,g10935);
  AN2 AND2_206(g28455,g27289,g20103);
  AN2 AND2_207(g33421,g32374,g21455);
  AN2 AND2_208(g21810,g3578,g20924);
  AN2 AND2_209(g17177,g6657,g14984);
  AN2 AND2_210(g21774,g3361,g20391);
  AN2 AND2_211(g29332,g29107,g22170);
  AN2 AND2_212(g23657,g19401,g11941);
  AN2 AND2_213(g28617,g27533,g20552);
  AN3 AND3_18(g34097,g33772,g9104,g18957);
  AN2 AND2_214(g21955,g5385,g21514);
  AN2 AND2_215(g23774,g14867,g21252);
  AN2 AND2_216(g22064,g15162,g19210);
  AN3 AND3_19(I24600,g6077,g6082,g9946);
  AN4 AND4_12(I31146,g30735,g31821,g32666,g32667);
  AN2 AND2_217(g25026,g22929,g10503);
  AN2 AND2_218(g34104,g33916,g23639);
  AN2 AND2_219(g27117,g26055,g16528);
  AN2 AND2_220(g21879,g4132,g19801);
  AN2 AND2_221(g34811,g14165,g34766);
  AN2 AND2_222(g21970,g5401,g21514);
  AN2 AND2_223(g18143,g586,g17533);
  AN2 AND2_224(g24502,g23428,g13223);
  AN2 AND2_225(g28201,g27499,g16720);
  AN2 AND2_226(g19536,g518,g16768);
  AN2 AND2_227(g19948,g17515,g16320);
  AN2 AND2_228(g29962,g23616,g28959);
  AN2 AND2_229(g21878,g4129,g19801);
  AN3 AND3_20(I16695,g10207,g12523,g12463);
  AN2 AND2_230(g32127,g31624,g29950);
  AN2 AND2_231(g31541,g22536,g29348);
  AN2 AND2_232(g24618,g22625,g19672);
  AN2 AND2_233(g26229,g1724,g25275);
  AN3 AND3_21(g33473,g32549,I31061,I31062);
  AN2 AND2_234(g18169,g676,g17433);
  AN2 AND2_235(g21886,g4153,g19801);
  AN2 AND2_236(g27568,g26576,g17791);
  AN2 AND2_237(g18791,g6044,g15634);
  AN2 AND2_238(g31789,g30201,g24013);
  AN2 AND2_239(g28467,g26993,g12295);
  AN2 AND2_240(g28494,g27973,g17741);
  AN2 AND2_241(g33789,g33159,g23022);
  AN2 AND2_242(g21792,g3396,g20391);
  AN2 AND2_243(g16591,g5256,g14879);
  AN2 AND2_244(g22009,g5782,g21562);
  AN2 AND2_245(g22665,g17174,g20905);
  AN2 AND2_246(g18168,g681,g17433);
  AN2 AND2_247(g18410,g2079,g15373);
  AN2 AND2_248(g21967,g5456,g21514);
  AN2 AND2_249(g21994,g5607,g19074);
  AN2 AND2_250(g31788,g21352,g29385);
  AN2 AND2_251(g33724,g14145,g33258);
  AN2 AND2_252(g32376,g2689,g31710);
  AN2 AND2_253(g19564,g17175,g13976);
  AN2 AND2_254(g33359,g32252,g20853);
  AN2 AND2_255(g25149,g14030,g23546);
  AN2 AND2_256(g17693,g1306,g13291);
  AN2 AND2_257(g22008,g5774,g21562);
  AN2 AND2_258(g32103,g31609,g29905);
  AN2 AND2_259(g24286,g4405,g22550);
  AN2 AND2_260(g18479,g2449,g15426);
  AN2 AND2_261(g18666,g4593,g17367);
  AN2 AND2_262(g33829,g33240,g20164);
  AN2 AND2_263(g18363,g1840,g17955);
  AN2 AND2_264(g32095,g7619,g30825);
  AN2 AND2_265(g18217,g15063,g16100);
  AN2 AND2_266(g33434,g32239,g29702);
  AN2 AND2_267(g24306,g4483,g22228);
  AN2 AND2_268(g33358,g32249,g20778);
  AN2 AND2_269(g25148,g16867,g23545);
  AN2 AND2_270(g11496,g4382,g7495);
  AN2 AND2_271(g15871,g3203,g13951);
  AN2 AND2_272(g18478,g2445,g15426);
  AN2 AND2_273(g30133,g28591,g21179);
  AN2 AND2_274(g33828,g33090,g24411);
  AN2 AND2_275(g28352,g10014,g27705);
  AN4 AND4_13(g11111,g5297,g7004,g5283,g9780);
  AN2 AND2_276(g14875,g1495,g10939);
  AN2 AND2_277(g34133,g33845,g23958);
  AN2 AND2_278(g21919,g15144,g21468);
  AN2 AND2_279(g30229,g28716,g23904);
  AN2 AND2_280(g25104,g16800,g23504);
  AN2 AND2_281(g11978,g2629,g7462);
  AN2 AND2_282(g26310,g2102,g25389);
  AN2 AND2_283(g23919,g4122,g19546);
  AN2 AND2_284(g32181,g31020,g19912);
  AN2 AND2_285(g33121,g8748,g32212);
  AN2 AND2_286(g18486,g2485,g15426);
  AN2 AND2_287(g27230,g25906,g19558);
  AN2 AND2_288(g27293,g9972,g26655);
  AN2 AND2_289(g29613,g28208,g19763);
  AN2 AND2_290(g28266,g23748,g27714);
  AN2 AND2_291(g19062,g446,g16180);
  AN2 AND2_292(g33344,g32228,g20670);
  AN2 AND2_293(g14218,g875,g10632);
  AN2 AND2_294(g21918,g5097,g21468);
  AN2 AND2_295(g30228,g28715,g23903);
  AN2 AND2_296(g26379,g19904,g25546);
  AN2 AND2_297(g18556,g2823,g15277);
  AN2 AND2_298(g25971,g1917,g24992);
  AN2 AND2_299(g24187,g305,g22722);
  AN2 AND2_300(g34228,g33750,g22942);
  AN2 AND2_301(g30011,g29183,g12930);
  AN2 AND2_302(g27265,g26785,g26759);
  AN4 AND4_14(I31226,g29385,g32781,g32782,g32783);
  AN2 AND2_303(g16844,g7212,g13000);
  AN2 AND2_304(g18580,g2907,g16349);
  AN2 AND2_305(g26050,g9630,g25047);
  AN4 AND4_15(g27416,g8046,g26314,g9187,g504);
  AN2 AND2_306(g26378,g19576,g25544);
  AN2 AND2_307(g13384,g4944,g11804);
  AN2 AND2_308(g29605,g2445,g28973);
  AN2 AND2_309(g18223,g1030,g16100);
  AN2 AND2_310(g23599,g19050,g9104);
  AN2 AND2_311(g27992,g26800,g23964);
  AN2 AND2_312(g22074,g6239,g19210);
  AN2 AND2_313(g27391,g26549,g17505);
  AN2 AND2_314(g24143,g17694,g21659);
  AN2 AND2_315(g25368,g6946,g22408);
  AN2 AND2_316(g27510,g26576,g17687);
  AN2 AND2_317(g34582,g7764,g34313);
  AN2 AND2_318(g32190,g142,g31233);
  AN2 AND2_319(g26096,g9733,g25268);
  AN2 AND2_320(g29951,g1874,g28786);
  AN2 AND2_321(g18110,g441,g17015);
  AN2 AND2_322(g34310,g14003,g34162);
  AN2 AND2_323(g25850,g3502,g24636);
  AN2 AND2_324(g15911,g3111,g13530);
  AN2 AND2_325(g28588,g27489,g20499);
  AN2 AND2_326(g28524,g6821,g27084);
  AN4 AND4_16(I31127,g32638,g32639,g32640,g32641);
  AN2 AND2_327(g18321,g1620,g17873);
  AN3 AND3_22(g24884,g3401,g23555,I24051);
  AN2 AND2_328(g30925,g29908,g23309);
  AN2 AND2_329(g21817,g3606,g20924);
  AN2 AND2_330(g11019,g5092,g9036);
  AN2 AND2_331(g18179,g763,g17328);
  AN2 AND2_332(g13019,g194,g11737);
  AN2 AND2_333(g18531,g2719,g15277);
  AN2 AND2_334(g30112,g28566,g20919);
  AN2 AND2_335(g28477,g27966,g17676);
  AN2 AND2_336(g33760,g33143,g20328);
  AN2 AND2_337(g24410,g3817,g23139);
  AN2 AND2_338(g32089,g27261,g31021);
  AN2 AND2_339(g25229,g7636,g22654);
  AN2 AND2_340(g30050,g22545,g28126);
  AN2 AND2_341(g29795,g28344,g23257);
  AN3 AND3_23(g34112,g22957,g9104,g33778);
  AN3 AND3_24(g11018,g7655,g7643,g7627);
  AN2 AND2_342(g18178,g758,g17328);
  AN2 AND2_343(g18740,g4572,g17384);
  AN2 AND2_344(g26857,g25062,g25049);
  AN2 AND2_345(g34050,g33772,g22942);
  AN2 AND2_346(g21977,g5535,g19074);
  AN2 AND2_347(g22092,g6419,g18833);
  AN2 AND2_348(g23532,g19400,g11852);
  AN2 AND2_349(g23901,g19606,g7963);
  AN2 AND2_350(g34378,g13095,g34053);
  AN2 AND2_351(g16025,g446,g14063);
  AN3 AND3_25(g33506,g32788,I31226,I31227);
  AN3 AND3_26(I24530,g9501,g9733,g5747);
  AN2 AND2_352(g32088,g27241,g31070);
  AN2 AND2_353(g24666,g11753,g22975);
  AN2 AND2_354(g22518,g12982,g19398);
  AN2 AND2_355(g21783,g3419,g20391);
  AN4 AND4_17(I31297,g32884,g32885,g32886,g32887);
  AN2 AND2_356(g24217,g18200,g22594);
  AN2 AND2_357(g18186,g753,g17328);
  AN2 AND2_358(g15785,g3558,g14107);
  AN2 AND2_359(g18676,g4358,g15758);
  AN2 AND2_360(g18685,g4688,g15885);
  AN2 AND2_361(g34386,g10800,g34060);
  AN2 AND2_362(g18373,g1890,g15171);
  AN2 AND2_363(g29514,g1608,g28780);
  AN2 AND2_364(g24015,g19540,g10951);
  AN2 AND2_365(g30096,g28546,g20770);
  AN2 AND2_366(g22637,g19363,g19489);
  AN2 AND2_367(g17176,g8616,g13008);
  AN2 AND2_368(g34742,g9000,g34698);
  AN2 AND2_369(g28616,g27532,g20551);
  AN3 AND3_27(g34096,g22957,g9104,g33772);
  AN2 AND2_370(g18654,g4146,g16249);
  AN2 AND2_371(g16203,g5821,g14297);
  AN2 AND2_372(g28313,g27231,g19766);
  AN2 AND2_373(g27116,g26026,g16527);
  AN4 AND4_18(I27509,g24084,g24085,g24086,g24087);
  AN2 AND2_374(g21823,g3731,g20453);
  AN2 AND2_375(g27615,g26789,g26770);
  AN2 AND2_376(g18800,g6187,g15348);
  AN2 AND2_377(g15859,g3610,g13923);
  AN4 AND4_19(I31181,g29385,g32716,g32717,g32718);
  AN2 AND2_378(g18417,g2116,g15373);
  AN2 AND2_379(g24556,g4035,g23341);
  AN2 AND2_380(g28285,g9657,g27717);
  AN2 AND2_381(g34681,g34491,g19438);
  AN4 AND4_20(I27508,g19935,g24082,g24083,g28033);
  AN2 AND2_382(g15858,g3542,g14045);
  AN2 AND2_383(g27041,g8519,g26330);
  AN2 AND2_384(g32126,g31601,g29948);
  AN2 AND2_385(g18334,g1696,g17873);
  AN2 AND2_386(g27275,g25945,g19745);
  AN2 AND2_387(g19756,g9899,g17154);
  AN2 AND2_388(g33927,g33094,g21412);
  AN3 AND3_28(g28254,g7268,g1668,g27395);
  AN2 AND2_389(g27430,g26488,g17579);
  AN2 AND2_390(g34857,g16540,g34813);
  AN2 AND2_391(g10822,g4264,g8514);
  AN2 AND2_392(g24223,g239,g22594);
  AN2 AND2_393(g27493,g246,g26837);
  AN2 AND2_394(g16957,g13064,g10418);
  AN2 AND2_395(g25959,g1648,g24963);
  AN2 AND2_396(g30730,g26346,g29778);
  AN2 AND2_397(g25925,g24990,g23234);
  AN2 AND2_398(g28466,g27960,g17637);
  AN2 AND2_399(g25112,g10428,g23510);
  AN2 AND2_400(g21966,g5406,g21514);
  AN2 AND2_401(g18762,g5475,g17929);
  AN2 AND2_402(g25050,g13056,g22312);
  AN2 AND2_403(g20084,g11591,g16609);
  AN2 AND2_404(g32339,g31474,g20672);
  AN2 AND2_405(g31240,g14793,g30206);
  AN2 AND2_406(g19350,g15968,g13505);
  AN2 AND2_407(g34765,g34692,g20057);
  AN2 AND2_408(g27340,g10199,g26784);
  AN2 AND2_409(g27035,g26348,g1500);
  AN2 AND2_410(g18423,g12851,g18008);
  AN2 AND2_411(g29789,g28270,g10233);
  AN2 AND2_412(g32338,g31466,g20668);
  AN3 AND3_29(g33491,g32679,I31151,I31152);
  AN2 AND2_413(g33903,g33447,g19146);
  AN2 AND2_414(g24922,g4831,g23931);
  AN2 AND2_415(g26129,g2384,g25121);
  AN2 AND2_416(g18216,g967,g15979);
  AN2 AND2_417(g24321,g4558,g22228);
  AN2 AND2_418(g16699,g7134,g12933);
  AN2 AND2_419(g27684,g26386,g20657);
  AN2 AND2_420(g28642,g27555,g20598);
  AN2 AND2_421(g18587,g2980,g16349);
  AN2 AND2_422(g25096,g23778,g20560);
  AN2 AND2_423(g29788,g28335,g23250);
  AN2 AND2_424(g26128,g2319,g25120);
  AN2 AND2_425(g14589,g10586,g10569);
  AN2 AND2_426(g29535,g2303,g28871);
  AN4 AND4_21(I31211,g31021,g31833,g32759,g32760);
  AN2 AND2_427(g27517,g26400,g17707);
  AN2 AND2_428(g10588,g7004,g5297);
  AN2 AND2_429(g18909,g16226,g13570);
  AN2 AND2_430(g32197,g31144,g20088);
  AN2 AND2_431(g18543,g2779,g15277);
  AN2 AND2_432(g26323,g10262,g25273);
  AN2 AND2_433(g24186,g18102,g22722);
  AN2 AND2_434(g14588,g11957,g11974);
  AN2 AND2_435(g24676,g2748,g23782);
  AN3 AND3_30(I16721,g10224,g12589,g12525);
  AN2 AND2_436(g18117,g464,g17015);
  AN2 AND2_437(g16427,g5216,g14876);
  AN2 AND2_438(g25802,g8106,g24586);
  AN2 AND2_439(g22083,g6287,g19210);
  AN2 AND2_440(g32411,g31119,g13469);
  AN2 AND2_441(g23023,g650,g20248);
  AN2 AND2_442(g19691,g9614,g17085);
  AN2 AND2_443(g24654,g11735,g22922);
  AN2 AND2_444(g28630,g27544,g20575);
  AN2 AND2_445(g29344,g29168,g18932);
  AN2 AND2_446(g18569,g94,g16349);
  AN2 AND2_447(g30002,g28481,g23487);
  AN2 AND2_448(g27130,g26026,g16585);
  AN2 AND2_449(g30057,g29144,g9462);
  AN2 AND2_450(g22622,g19336,g19469);
  AN2 AND2_451(g18568,g37,g16349);
  AN2 AND2_452(g18747,g5138,g17847);
  AN2 AND2_453(g25765,g24989,g24973);
  AN2 AND2_454(g27362,g26080,g20036);
  AN2 AND2_455(g31990,g31772,g18945);
  AN2 AND2_456(g33899,g32132,g33335);
  AN2 AND2_457(g18242,g962,g16431);
  AN2 AND2_458(g10616,g7998,g174);
  AN2 AND2_459(g27523,g26549,g17718);
  AN2 AND2_460(g30245,g28733,g23935);
  AN4 AND4_22(I31126,g30673,g31818,g32636,g32637);
  AN2 AND2_461(g26232,g2193,g25396);
  AN2 AND2_462(g33898,g33419,g15655);
  AN2 AND2_463(g21816,g3602,g20924);
  AN2 AND2_464(g18123,g479,g16886);
  AN2 AND2_465(g18814,g6519,g15483);
  AN2 AND2_466(g33719,g33141,g19433);
  AN2 AND2_467(g24762,g655,g23573);
  AN3 AND3_31(g10704,g2145,g10200,g2130);
  AN2 AND2_468(g34533,g34318,g19731);
  AN2 AND2_469(g18751,g5156,g17847);
  AN2 AND2_470(g18807,g6386,g15656);
  AN2 AND2_471(g21976,g5527,g19074);
  AN2 AND2_472(g21985,g5571,g19074);
  AN2 AND2_473(g15902,g441,g13975);
  AN2 AND2_474(g18772,g5689,g15615);
  AN2 AND2_475(g28555,g27429,g20373);
  AN2 AND2_476(g33718,g33147,g19432);
  AN2 AND2_477(g34298,g8679,g34132);
  AN2 AND2_478(g28454,g26976,g12233);
  AN3 AND3_32(g33521,g32895,I31301,I31302);
  AN2 AND2_479(g18974,g174,g16127);
  AN4 AND4_23(g26261,g24688,g10678,g8778,g8757);
  AN2 AND2_480(g32315,g31306,g23517);
  AN2 AND2_481(g24423,g4950,g22897);
  AN2 AND2_482(g21752,g3171,g20785);
  AN4 AND4_24(g27727,g22432,g25211,g26424,g26195);
  AN4 AND4_25(I31296,g30937,g31848,g32882,g32883);
  AN2 AND2_483(g18639,g3831,g17096);
  AN2 AND2_484(g28570,g27456,g20434);
  AN2 AND2_485(g28712,g27590,g20708);
  AN2 AND2_486(g21954,g5381,g21514);
  AN2 AND2_487(g27222,g26055,g13932);
  AN2 AND2_488(g29760,g28309,g23227);
  AN2 AND2_489(g33832,g33088,g27991);
  AN2 AND2_490(g18230,g1111,g16326);
  AN4 AND4_26(g29029,g14506,g25227,g26424,g27494);
  AN2 AND2_491(g17139,g8635,g12967);
  AN2 AND2_492(g18293,g1484,g16449);
  AN4 AND4_27(g17653,g11547,g11592,g6789,I18620);
  AN2 AND2_493(g15738,g1111,g13260);
  AN2 AND2_494(g18638,g3827,g17096);
  AN2 AND2_495(g27437,g26576,g17589);
  AN2 AND2_496(g33440,g32250,g29719);
  AN2 AND2_497(g32055,g10999,g30825);
  AN2 AND2_498(g17138,g255,g13239);
  AN2 AND2_499(g18265,g1270,g16000);
  AN2 AND2_500(g25129,g17682,g23527);
  AN2 AND2_501(g15699,g1437,g13861);
  AN2 AND2_502(g30232,g28719,g23912);
  AN2 AND2_503(g32111,g31616,g29922);
  AN2 AND2_504(g18416,g2112,g15373);
  AN2 AND2_505(g25057,g23275,g20511);
  AN2 AND2_506(g32070,g10967,g30825);
  AN2 AND2_507(g33861,g33271,g20502);
  AN2 AND2_508(g28239,g27135,g19659);
  AN2 AND2_509(g25128,g17418,g23525);
  AN2 AND2_510(g17636,g10829,g13463);
  AN2 AND2_511(g11916,g2227,g7328);
  AN2 AND2_512(g33247,g32130,g19980);
  AN2 AND2_513(g28567,g6832,g27101);
  AN4 AND4_28(I31197,g32740,g32741,g32742,g32743);
  AN2 AND2_514(g27347,g26400,g17390);
  AN2 AND2_515(g18992,g8341,g16171);
  AN2 AND2_516(g18391,g1982,g15171);
  AN3 AND3_33(g24908,g3752,g23239,I24075);
  AN2 AND2_517(g28238,g27133,g19658);
  AN2 AND2_518(g21842,g3863,g21070);
  AN2 AND2_519(g18510,g2625,g15509);
  AN2 AND2_520(g30261,g28772,g23961);
  AN2 AND2_521(g23392,g7247,g21430);
  AN2 AND2_522(g24569,g5115,g23382);
  AN2 AND2_523(g25323,g6888,g22359);
  AN2 AND2_524(g31324,g30171,g27937);
  AN2 AND2_525(g33099,g32395,g18944);
  AN2 AND2_526(g13287,g1221,g11472);
  AN2 AND2_527(g27600,g26755,g26725);
  AN4 AND4_29(g10733,g3639,g6905,g3625,g8542);
  AN2 AND2_528(g18579,g2984,g16349);
  AN2 AND2_529(g31777,g21343,g29385);
  AN2 AND2_530(g33701,g33162,g16305);
  AN2 AND2_531(g24747,g17510,g22417);
  AN2 AND2_532(g32067,g4727,g30614);
  AN2 AND2_533(g21559,g16236,g10897);
  AN2 AND2_534(g31272,g30117,g27742);
  AN3 AND3_34(I16618,g10124,g12341,g12293);
  AN2 AND2_535(g15632,g3494,g13555);
  AN2 AND2_536(g28185,g27026,g19435);
  AN3 AND3_35(g10874,g7791,g6219,g6227);
  AN2 AND2_537(g18578,g2873,g16349);
  AN2 AND2_538(g25775,g2922,g24568);
  AN2 AND2_539(g23424,g7345,g21556);
  AN2 AND2_540(g27351,g10218,g26804);
  AN2 AND2_541(g27372,g26488,g17476);
  AN2 AND2_542(g19768,g2803,g15833);
  AN2 AND2_543(g14874,g1099,g10909);
  AN2 AND2_544(g16671,g6275,g14817);
  AN2 AND2_545(g21558,g15904,g13729);
  AN2 AND2_546(g27821,g7680,g25892);
  AN2 AND2_547(g32150,g31624,g29995);
  AN2 AND2_548(g28154,g8492,g27306);
  AN2 AND2_549(g18586,g2886,g16349);
  AN2 AND2_550(g29649,g2241,g28678);
  AN3 AND3_36(g33462,g32470,I31006,I31007);
  AN2 AND2_551(g21830,g3774,g20453);
  AN2 AND2_552(g26611,g24935,g20580);
  AN2 AND2_553(g20751,g16260,g4836);
  AN2 AND2_554(g10665,g209,g8292);
  AN2 AND2_555(g28637,g22399,g27011);
  AN2 AND2_556(g18442,g2259,g18008);
  AN2 AND2_557(g32019,g30579,g22358);
  AN2 AND2_558(g24772,g16287,g23061);
  AN2 AND2_559(g29648,g2112,g29121);
  AN2 AND2_560(g27264,g25941,g19714);
  AN2 AND2_561(g22115,g6573,g19277);
  AN2 AND2_562(g27137,g26026,g16606);
  AN2 AND2_563(g21865,g3965,g21070);
  AN2 AND2_564(g31140,g2102,g30037);
  AN2 AND2_565(g32196,g27587,g31376);
  AN2 AND2_566(g13942,g5897,g12512);
  AN2 AND2_567(g24639,g6181,g23699);
  AN2 AND2_568(g32018,g4146,g30937);
  AN2 AND2_569(g26271,g1992,g25341);
  AN2 AND2_570(g29604,g2315,g28966);
  AN3 AND3_37(g30316,g29199,g7097,g6682);
  AN2 AND2_571(g21713,g298,g20283);
  AN2 AND2_572(g34499,g31288,g34339);
  AN2 AND2_573(g24230,g901,g22594);
  AN3 AND3_38(g13156,g10816,g10812,g10805);
  AN2 AND2_574(g18116,g168,g17015);
  AN2 AND2_575(g24293,g4438,g22550);
  AN2 AND2_576(g18615,g3347,g17200);
  AN2 AND2_577(g22052,g6113,g21611);
  AN3 AND3_39(g10476,g7244,g7259,I13862);
  AN2 AND2_578(g24638,g22763,g19690);
  AN2 AND2_579(g29770,g28320,g23238);
  AN2 AND2_580(g16190,g14626,g11810);
  AN2 AND2_581(g29563,g1616,g28853);
  AN4 AND4_30(I31202,g32747,g32748,g32749,g32750);
  AN2 AND2_582(g34498,g13888,g34336);
  AN2 AND2_583(g18720,g15137,g16795);
  AN2 AND2_584(g26753,g16024,g24452);
  AN4 AND4_31(I31257,g32826,g32827,g32828,g32829);
  AN2 AND2_585(g25880,g8443,g24814);
  AN4 AND4_32(g14555,g12521,g12356,g12307,I16671);
  AN2 AND2_586(g24416,g4939,g22870);
  AN2 AND2_587(g16520,g5909,g14965);
  AN2 AND2_588(g21705,g209,g20283);
  AN2 AND2_589(g30056,g29165,g12659);
  AN2 AND2_590(g18275,g15070,g16136);
  AN2 AND2_591(g26145,g11962,g25131);
  AN4 AND4_33(I31111,g31070,g31815,g32615,g32616);
  AN2 AND2_592(g18430,g2204,g18008);
  AN2 AND2_593(g18746,g5134,g17847);
  AN3 AND3_40(g27209,g26213,g8365,g2051);
  AN2 AND2_594(g32402,g4888,g30990);
  AN2 AND2_595(g18493,g2514,g15426);
  AN2 AND2_596(g33871,g33281,g20546);
  AN2 AND2_597(g30080,g28121,g20674);
  AN2 AND2_598(g28215,g9264,g27565);
  AN2 AND2_599(g26650,g10796,g24424);
  AN3 AND3_41(g34080,g22957,g9104,g33750);
  AN2 AND2_600(g16211,g5445,g14215);
  AN2 AND2_601(g27208,g9037,g26598);
  AN2 AND2_602(g18465,g2384,g15224);
  AN2 AND2_603(g29767,g28317,g23236);
  AN2 AND2_604(g29794,g28342,g23256);
  AN2 AND2_605(g21188,g7666,g15705);
  AN2 AND2_606(g33360,g32253,g20869);
  AN2 AND2_607(g18237,g1146,g16326);
  AN2 AND2_608(g29845,g28375,g23291);
  AN2 AND2_609(g23188,g13994,g20025);
  AN3 AND3_42(I16143,g8751,g11491,g11445);
  AN2 AND2_610(g28439,g27273,g10233);
  AN2 AND2_611(g18340,g1720,g17873);
  AN2 AND2_612(g29899,g28428,g23375);
  AN2 AND2_613(g29990,g29007,g9239);
  AN2 AND2_614(g21939,g5224,g18997);
  AN2 AND2_615(g25831,g3151,g24623);
  AN2 AND2_616(g15784,g3235,g13977);
  AN2 AND2_617(g18806,g6381,g15656);
  AN2 AND2_618(g18684,g4681,g15885);
  AN2 AND2_619(g26393,g19467,g25558);
  AN2 AND2_620(g14567,g10568,g10552);
  AN2 AND2_621(g24835,g8720,g23233);
  AN2 AND2_622(g29633,g1978,g29085);
  AN4 AND4_34(I31067,g32552,g32553,g32554,g32555);
  AN2 AND2_623(g24014,g7933,g19063);
  AN2 AND2_624(g15103,g4180,g14454);
  AN2 AND2_625(g34753,g34676,g19586);
  AN2 AND2_626(g21938,g5216,g18997);
  AN2 AND2_627(g18142,g577,g17533);
  AN2 AND2_628(g34342,g34103,g19998);
  AN2 AND2_629(g30145,g28603,g21247);
  AN2 AND2_630(g30031,g29071,g10540);
  AN2 AND2_631(g27614,g26785,g26759);
  AN2 AND2_632(g32256,g31249,g20382);
  AN2 AND2_633(g18517,g2652,g15509);
  AN2 AND2_634(g27436,g26576,g17588);
  AN2 AND2_635(g30199,g28664,g23861);
  AN2 AND2_636(g29718,g28512,g11136);
  AN2 AND2_637(g29521,g1744,g28824);
  AN2 AND2_638(g16700,g5208,g14838);
  AN2 AND2_639(g31220,g30273,g25202);
  AN3 AND3_43(g33472,g32542,I31056,I31057);
  AN2 AND2_640(g16126,g5495,g14262);
  AN2 AND2_641(g28284,g11398,g27994);
  AN2 AND2_642(g10675,g3436,g8500);
  AN2 AND2_643(g25989,g25258,g21012);
  AN4 AND4_35(g27073,g7121,g3873,g3881,g26281);
  AN2 AND2_644(g30198,g28662,g23860);
  AN2 AND2_645(g32300,g31274,g20544);
  AN2 AND2_646(g14185,g8686,g11744);
  AN2 AND2_647(g25056,g12779,g23456);
  AN2 AND2_648(g28304,g27226,g19753);
  AN2 AND2_649(g33911,g33137,g10725);
  AN2 AND2_650(g34198,g33688,g24491);
  AN2 AND2_651(g26161,g2518,g25139);
  AN2 AND2_652(g34529,g34306,g19634);
  AN2 AND2_653(g21875,g4116,g19801);
  AN2 AND2_654(g25988,g9510,g25016);
  AN4 AND4_36(I31196,g30825,g31830,g32738,g32739);
  AN2 AND2_655(g25924,g24976,g16846);
  AN2 AND2_656(g27346,g26400,g17389);
  AN2 AND2_657(g34528,g34305,g19617);
  AN2 AND2_658(g17692,g1124,g13307);
  AN2 AND2_659(g18130,g528,g16971);
  AN2 AND2_660(g34696,g34531,g20004);
  AN2 AND2_661(g18193,g837,g17821);
  AN2 AND2_662(g22013,g5802,g21562);
  AN2 AND2_663(g32157,g31646,g30021);
  AN2 AND2_664(g34393,g34189,g21304);
  AN2 AND2_665(g26259,g24430,g25232);
  AN3 AND3_44(I24508,g9434,g9672,g5401);
  AN2 AND2_666(g18362,g1834,g17955);
  AN2 AND2_667(g23218,g20200,g16530);
  AN2 AND2_668(g29861,g28390,g23313);
  AN2 AND2_669(g29573,g1752,g28892);
  AN2 AND2_670(g33071,g31591,g32404);
  AN2 AND2_671(g21837,g3719,g20453);
  AN2 AND2_672(g34764,g34691,g20009);
  AN2 AND2_673(g22329,g11940,g20329);
  AN2 AND2_674(g10883,g3355,g9061);
  AN2 AND2_675(g18165,g650,g17433);
  AN2 AND2_676(g23837,g21160,g10804);
  AN2 AND2_677(g18523,g2675,g15509);
  AN2 AND2_678(g26087,g5475,g25072);
  AN2 AND2_679(g27034,g26328,g8609);
  AN2 AND2_680(g13306,g441,g11048);
  AN2 AND2_681(g31776,g21329,g29385);
  AN2 AND2_682(g34365,g34149,g20451);
  AN2 AND2_683(g26258,g12875,g25231);
  AN2 AND2_684(g19651,g1111,g16119);
  AN2 AND2_685(g33785,g33100,g20550);
  AN2 AND2_686(g29926,g1604,g28736);
  AN2 AND2_687(g34869,g34816,g19869);
  AN2 AND2_688(g28139,g27337,g26054);
  AN2 AND2_689(g22005,g5759,g21562);
  AN2 AND2_690(g31147,g12286,g30054);
  AN2 AND2_691(g28653,g7544,g27014);
  AN2 AND2_692(g13038,g8509,g11034);
  AN2 AND2_693(g27292,g1714,g26654);
  AN2 AND2_694(g29612,g27875,g28633);
  AN2 AND2_695(g24465,g3827,g23139);
  AN3 AND3_45(g12641,g10295,g3171,g3179);
  AN2 AND2_696(g22538,g14035,g20248);
  AN2 AND2_697(g27153,g26055,g16629);
  AN2 AND2_698(g33355,g32243,g20769);
  AN2 AND2_699(g29324,g29078,g18883);
  AN2 AND2_700(g34868,g34813,g19866);
  AN2 AND2_701(g7396,g392,g441);
  AN2 AND2_702(g25031,g20675,g23432);
  AN2 AND2_703(g30161,g28614,g21275);
  AN2 AND2_704(g18475,g12853,g15426);
  AN2 AND2_705(g33859,g33426,g10531);
  AN4 AND4_37(g26244,g24688,g8812,g10658,g8757);
  AN2 AND2_706(g29534,g28965,g22457);
  AN2 AND2_707(g33370,g32279,g21139);
  AN2 AND2_708(g24983,g23217,g20238);
  AN2 AND2_709(g27409,g26519,g17524);
  AN2 AND2_710(g16855,g4392,g13107);
  AN2 AND2_711(g18727,g4931,g16077);
  AN2 AND2_712(g28415,g27250,g19963);
  AN2 AND2_713(g24684,g11769,g22989);
  AN2 AND2_714(g28333,g27239,g19787);
  AN2 AND2_715(g33858,g33268,g20448);
  AN2 AND2_716(g34709,g34549,g17242);
  AN2 AND2_717(g18222,g1024,g16100);
  AN2 AND2_718(g10501,g1233,g9007);
  AN2 AND2_719(g16870,g6625,g14905);
  AN2 AND2_720(g27136,g26026,g16605);
  AN2 AND2_721(g27408,g26519,g17523);
  AN4 AND4_38(g27635,g23032,g26281,g26424,g24996);
  AN2 AND2_722(g21915,g5080,g21468);
  AN2 AND2_723(g30225,g28705,g23897);
  AN2 AND2_724(g31151,g10037,g30065);
  AN2 AND2_725(g18437,g2241,g18008);
  AN2 AND2_726(g24142,g17700,g21657);
  AN4 AND4_39(I31001,g29385,g32456,g32457,g32458);
  AN2 AND2_727(g31996,g31779,g18979);
  AN2 AND2_728(g34225,g33744,g22942);
  AN4 AND4_40(I31077,g32566,g32567,g32568,g32569);
  AN2 AND2_729(g26602,g7487,g24453);
  AN2 AND2_730(g30258,g28751,g23953);
  AN2 AND2_731(g11937,g1936,g7362);
  AN2 AND2_732(g15860,g3889,g14160);
  AN3 AND3_46(g34087,g33766,g9104,g18957);
  AN2 AND2_733(g23201,g14027,g20040);
  AN2 AND2_734(g33844,g33257,g20327);
  AN2 AND2_735(g33367,g32271,g21053);
  AN4 AND4_41(I31256,g31021,g31841,g32824,g32825);
  AN2 AND2_736(g18703,g4776,g16782);
  AN2 AND2_737(g22100,g6466,g18833);
  AN2 AND2_738(g18347,g1756,g17955);
  AN2 AND2_739(g19717,g6527,g17122);
  AN2 AND2_740(g14438,g1087,g10726);
  AN2 AND2_741(g30043,g29106,g9392);
  AN2 AND2_742(g18253,g1211,g16897);
  AN2 AND2_743(g25132,g10497,g23528);
  AN2 AND2_744(g30244,g28732,g23930);
  AN4 AND4_42(g26171,g25357,g6856,g11709,g11686);
  AN2 AND2_745(g15700,g3089,g13483);
  AN3 AND3_47(I24051,g3380,g3385,g8492);
  AN2 AND2_746(g18600,g3111,g16987);
  AN2 AND2_747(g20193,g15578,g17264);
  AN2 AND2_748(g18781,g5831,g18065);
  AN2 AND2_749(g28585,g27063,g10530);
  AN2 AND2_750(g24193,g336,g22722);
  AN4 AND4_43(g28484,g27187,g10290,g21163,I26972);
  AN2 AND2_751(g33420,g32373,g21454);
  AN2 AND2_752(g30069,g29175,g12708);
  AN2 AND2_753(g29766,g28316,g23235);
  AN2 AND2_754(g18236,g15065,g16326);
  AN2 AND2_755(g21782,g3416,g20391);
  AN2 AND2_756(g17771,g13288,g13190);
  AN2 AND2_757(g20165,g5156,g17733);
  AN2 AND2_758(g34069,g8774,g33797);
  AN2 AND2_759(g21984,g5563,g19074);
  AN4 AND4_44(I31102,g32603,g32604,g32605,g32606);
  AN4 AND4_45(g26994,g23032,g26226,g26424,g25557);
  AN4 AND4_46(g27474,g8038,g26314,g518,g504);
  AN2 AND2_760(g28554,g27426,g20372);
  AN4 AND4_47(I31157,g32682,g32683,g32684,g32685);
  AN2 AND2_761(g18351,g1760,g17955);
  AN2 AND2_762(g18372,g1886,g15171);
  AN2 AND2_763(g24523,g22318,g19468);
  AN2 AND2_764(g32314,g31304,g23516);
  AN2 AND2_765(g29871,g28400,g23332);
  AN2 AND2_766(g33446,g32385,g21607);
  AN4 AND4_48(g27711,g22369,g25193,g26424,g26166);
  AN2 AND2_767(g16707,g6641,g15033);
  AN2 AND2_768(g21419,g16681,g13595);
  AN2 AND2_769(g32287,g2823,g30578);
  AN2 AND2_770(g34774,g34695,g20180);
  AN2 AND2_771(g18175,g744,g17328);
  AN2 AND2_772(g18821,g15168,g15680);
  AN2 AND2_773(g34955,g34931,g34320);
  AN2 AND2_774(g27327,g2116,g26732);
  AN2 AND2_775(g34375,g13077,g34049);
  AN2 AND2_776(g16202,g86,g14197);
  AN2 AND2_777(g28312,g27828,g26608);
  AN2 AND2_778(g28200,g27652,g11383);
  AN2 AND2_779(g32307,g31291,g23500);
  AN2 AND2_780(g14566,g10566,g10551);
  AN2 AND2_781(g32085,g27253,g31021);
  AN4 AND4_49(I31066,g31070,g31807,g32550,g32551);
  AN2 AND2_782(g29360,g27364,g28294);
  AN2 AND2_783(g21822,g3727,g20453);
  AN2 AND2_784(g22515,g12981,g19395);
  AN4 AND4_50(I31231,g31376,g31836,g32789,g32790);
  AN2 AND2_785(g22991,g645,g20248);
  AN2 AND2_786(g27537,g26549,g17742);
  AN2 AND2_787(g28115,g27354,g22759);
  AN2 AND2_788(g31540,g29904,g23548);
  AN2 AND2_789(g25087,g17307,g23489);
  AN2 AND2_790(g32054,g10890,g30735);
  AN2 AND2_791(g24475,g3831,g23139);
  AN2 AND2_792(g7685,g4382,g4375);
  AN2 AND2_793(g18264,g1263,g16000);
  AN2 AND2_794(g18790,g6040,g15634);
  AN2 AND2_795(g18137,g538,g17249);
  AN4 AND4_51(I27513,g19984,g24089,g24090,g28034);
  AN2 AND2_796(g18516,g2638,g15509);
  AN2 AND2_797(g34337,g34095,g19881);
  AN2 AND2_798(g24727,g13300,g23016);
  AN2 AND2_799(g34171,g33925,g24360);
  AN2 AND2_800(g16590,g5236,g14683);
  AN2 AND2_801(g24222,g262,g22594);
  AN2 AND2_802(g16986,g246,g13142);
  AN2 AND2_803(g27303,g11996,g26681);
  AN2 AND2_804(g11223,g8281,g8505);
  AN2 AND2_805(g25043,g20733,g23447);
  AN2 AND2_806(g32269,g31253,g20443);
  AN2 AND2_807(g21853,g3917,g21070);
  AN4 AND4_52(g28799,g21434,g26424,g25348,g27445);
  AN2 AND2_808(g26079,g6199,g25060);
  AN2 AND2_809(g34967,g34951,g23189);
  AN2 AND2_810(g28813,g4104,g27038);
  AN2 AND2_811(g29629,g28211,g19779);
  AN2 AND2_812(g32341,g31472,g23610);
  AN2 AND2_813(g31281,g30106,g27742);
  AN2 AND2_814(g15870,g3231,g13948);
  AN2 AND2_815(g26078,g5128,g25055);
  AN2 AND2_816(g32156,g31639,g30018);
  AN2 AND2_817(g25069,g23296,g20535);
  AN2 AND2_818(g24703,g17592,g22369);
  AN2 AND2_819(g31301,g30170,g27907);
  AN2 AND2_820(g18209,g921,g15938);
  AN2 AND2_821(g29628,g27924,g28648);
  AN2 AND2_822(g33902,g33085,g13202);
  AN2 AND2_823(g21836,g3805,g20453);
  AN2 AND2_824(g31120,g1700,g29976);
  AN2 AND2_825(g32180,g2791,g31638);
  AN2 AND2_826(g23836,g4129,g19495);
  AN2 AND2_827(g26086,g9672,g25255);
  AN2 AND2_828(g28674,g27569,g20629);
  AN2 AND2_829(g13321,g847,g11048);
  AN2 AND2_830(g25068,g17574,g23477);
  AN2 AND2_831(g25955,g24720,g19580);
  AN2 AND2_832(g30919,g29898,g23286);
  AN2 AND2_833(g18208,g930,g15938);
  AN2 AND2_834(g16801,g5120,g14238);
  AN2 AND2_835(g16735,g6235,g15027);
  AN2 AND2_836(g23401,g7262,g21460);
  AN2 AND2_837(g25879,g11135,g24683);
  AN2 AND2_838(g24600,g22591,g19652);
  AN2 AND2_839(g25970,g1792,g24991);
  AN2 AND2_840(g31146,g12285,g30053);
  AN2 AND2_841(g30010,g29035,g9274);
  AN2 AND2_842(g30918,g8681,g29707);
  AN2 AND2_843(g32335,g6199,g31566);
  AN4 AND4_53(g11178,g6682,g7097,g6668,g10061);
  AN2 AND2_844(g11740,g8769,g703);
  AN2 AND2_845(g18542,g2787,g15277);
  AN3 AND3_48(I18803,g13156,g11450,g6756);
  AN2 AND2_846(g18453,g2315,g15224);
  AN2 AND2_847(g29591,g28552,g11346);
  AN2 AND2_848(g29785,g28332,g23248);
  AN2 AND2_849(g31290,g29734,g23335);
  AN2 AND2_850(g22114,g6565,g19277);
  AN2 AND2_851(g26159,g2370,g25137);
  AN2 AND2_852(g26125,g1894,g25117);
  AN2 AND2_853(g21864,g3961,g21070);
  AN2 AND2_854(g34079,g33703,g19532);
  AN2 AND2_855(g22082,g6283,g19210);
  AN2 AND2_856(g27390,g26549,g17504);
  AN2 AND2_857(g18726,g4927,g16077);
  AN4 AND4_54(g26977,g23032,g26261,g26424,g25550);
  AN2 AND2_858(g30599,g18911,g29863);
  AN2 AND2_859(g22107,g6411,g18833);
  AN2 AND2_860(g30078,g28526,g20667);
  AN2 AND2_861(g21749,g3155,g20785);
  AN2 AND2_862(g26158,g2255,g25432);
  AN4 AND4_55(g17725,g11547,g11592,g6789,I18716);
  AN2 AND2_863(g26783,g25037,g21048);
  AN4 AND4_56(I31287,g32870,g32871,g32872,g32873);
  AN2 AND2_864(g18614,g3343,g17200);
  AN2 AND2_865(g28692,g27578,g20661);
  AN4 AND4_57(g28761,g21434,g26424,g25299,g27416);
  AN2 AND2_866(g34078,g33699,g19531);
  AN2 AND2_867(g18436,g2227,g18008);
  AN2 AND2_868(g25967,g9373,g24986);
  AN2 AND2_869(g30598,g18898,g29862);
  AN2 AND2_870(g14585,g1141,g10905);
  AN2 AND2_871(g29859,g28388,g23307);
  AN4 AND4_58(I31307,g32898,g32899,g32900,g32901);
  AN4 AND4_59(I31076,g30614,g31809,g32564,g32565);
  AN2 AND2_872(g30086,g28536,g20704);
  AN2 AND2_873(g21748,g15089,g20785);
  AN2 AND2_874(g15707,g4082,g13506);
  AN2 AND2_875(g15819,g3251,g14101);
  AN2 AND2_876(g18607,g3139,g16987);
  AN3 AND3_49(g34086,g20114,g33766,g9104);
  AN2 AND2_877(g18320,g1616,g17873);
  AN2 AND2_878(g24790,g7074,g23681);
  AN2 AND2_879(g21276,g10157,g17625);
  AN2 AND2_880(g21285,g7857,g16027);
  AN2 AND2_881(g26295,g13070,g25266);
  AN2 AND2_882(g29858,g28387,g23306);
  AN2 AND2_883(g21704,g164,g20283);
  AN2 AND2_884(g18274,g1311,g16031);
  AN2 AND2_885(g22849,g1227,g19653);
  AN2 AND2_886(g33366,g32268,g21010);
  AN2 AND2_887(g27522,g26549,g17717);
  AN2 AND2_888(g26823,g24401,g13106);
  AN2 AND2_889(g15818,g3941,g14082);
  AN2 AND2_890(g18530,g2715,g15277);
  AN3 AND3_50(g25459,g6058,g23844,I24582);
  AN2 AND2_891(g18593,g2999,g16349);
  AN2 AND2_892(g18346,g1752,g17955);
  AN2 AND2_893(g19716,g12100,g17121);
  AN2 AND2_894(g21809,g3574,g20924);
  AN2 AND2_895(g23254,g20056,g20110);
  AN2 AND2_896(g28214,g27731,g26625);
  AN2 AND2_897(g15111,g4281,g14454);
  AN2 AND2_898(g22848,g19449,g19649);
  AN2 AND2_899(g18122,g15052,g17015);
  AN2 AND2_900(g23900,g1129,g19408);
  AN2 AND2_901(g34322,g14188,g34174);
  AN4 AND4_60(g14608,g12638,g12476,g12429,I16721);
  AN2 AND2_902(g15978,g246,g14032);
  AN2 AND2_903(g18565,g2852,g16349);
  AN2 AND2_904(g26336,g10307,g25480);
  AN2 AND2_905(g30125,g28581,g21056);
  AN2 AND2_906(g18464,g2370,g15224);
  AN2 AND2_907(g21808,g3570,g20924);
  AN2 AND2_908(g29844,g28374,g23290);
  AN2 AND2_909(g34532,g34314,g19710);
  AN2 AND2_910(g15590,g3139,g13530);
  AN2 AND2_911(g29367,g8575,g28325);
  AN2 AND2_912(g28539,g27187,g12762);
  AN2 AND2_913(g10921,g1548,g8685);
  AN2 AND2_914(g27483,g26488,g17642);
  AN2 AND2_915(g30158,g28613,g21274);
  AN2 AND2_916(g33403,g32352,g21396);
  AN2 AND2_917(g24422,g4771,g22896);
  AN4 AND4_61(I31341,g31710,g31856,g32947,g32948);
  AN2 AND2_918(g32278,g2811,g30572);
  AN2 AND2_919(g27553,g26293,g23353);
  AN2 AND2_920(g18641,g3841,g17096);
  AN2 AND2_921(g18797,g6173,g15348);
  AN2 AND2_922(g25079,g21011,g23483);
  AN4 AND4_62(I31156,g31070,g31823,g32680,g32681);
  AN2 AND2_923(g18292,g1472,g16449);
  AN2 AND2_924(g16706,g6621,g14868);
  AN2 AND2_925(g31226,g30282,g25218);
  AN2 AND2_926(g32286,g31658,g29312);
  AN2 AND2_927(g34561,g34368,g17410);
  AN2 AND2_928(g16597,g6263,g15021);
  AN2 AND2_929(g18153,g626,g17533);
  AN2 AND2_930(g27326,g12048,g26731);
  AN2 AND2_931(g25078,g23298,g20538);
  AN2 AND2_932(g31481,g29768,g23417);
  AN2 AND2_933(g32039,g31476,g20070);
  AN2 AND2_934(g33715,g33135,g19416);
  AN2 AND2_935(g32306,g31289,g23499);
  AN2 AND2_936(g34295,g34057,g19370);
  AN3 AND3_51(g33481,g32607,I31101,I31102);
  AN2 AND2_937(g22135,g6657,g19277);
  AN2 AND2_938(g27536,g26519,g17738);
  AN2 AND2_939(g18409,g2084,g15373);
  AN4 AND4_63(g27040,g7812,g6565,g6573,g26226);
  AN2 AND2_940(g25086,g13941,g23488);
  AN2 AND2_941(g21733,g3034,g20330);
  AN3 AND3_52(g10674,g6841,g10200,g2130);
  AN2 AND2_942(g18136,g550,g17249);
  AN2 AND2_943(g18408,g2070,g15373);
  AN2 AND2_944(g18635,g3808,g17096);
  AN2 AND2_945(g24726,g15965,g23015);
  AN2 AND2_946(g27252,g26733,g26703);
  AN2 AND2_947(g24913,g4821,g23908);
  AN2 AND2_948(g21874,g4112,g19801);
  AN2 AND2_949(g25817,g24807,g21163);
  AN2 AND2_950(g32187,g30672,g25287);
  AN2 AND2_951(g26289,g2551,g25400);
  AN2 AND2_952(g24436,g3125,g23067);
  AN2 AND2_953(g25159,g4907,g22908);
  AN3 AND3_53(g10732,g6850,g2697,g2689);
  AN2 AND2_954(g22049,g6082,g21611);
  AN2 AND2_955(g25125,g20187,g23520);
  AN2 AND2_956(g27564,g26305,g23378);
  AN2 AND2_957(g25901,g24853,g16290);
  AN2 AND2_958(g26023,g9528,g25036);
  AN4 AND4_64(I31131,g31542,g31819,g32643,g32644);
  AN2 AND2_959(g34966,g34950,g23170);
  AN2 AND2_960(g31490,g29786,g23429);
  AN2 AND2_961(g10934,g9197,g7918);
  AN2 AND2_962(g24607,g5817,g23666);
  AN2 AND2_963(g25977,g25236,g20875);
  AN2 AND2_964(g26288,g2259,g25309);
  AN3 AND3_54(g33490,g32672,I31146,I31147);
  AN2 AND2_965(g19681,g5835,g17014);
  AN2 AND2_966(g24320,g6973,g22228);
  AN2 AND2_967(g28235,g9467,g27592);
  AN2 AND2_968(g26571,g10472,g24386);
  AN2 AND2_969(g23166,g13959,g19979);
  AN2 AND2_970(g23009,g20196,g14219);
  AN2 AND2_971(g22048,g6052,g21611);
  AN2 AND2_972(g26308,g6961,g25289);
  AN3 AND3_55(g29203,g24095,I27513,I27514);
  AN2 AND2_973(g18164,g699,g17433);
  AN2 AND2_974(g28683,g27876,g20649);
  AN2 AND2_975(g32143,g31646,g29967);
  AN2 AND2_976(g31784,g30176,g24003);
  AN2 AND2_977(g34364,g34048,g24366);
  AN2 AND2_978(g33784,g33107,g20531);
  AN2 AND2_979(g31376,g24952,g29814);
  AN2 AND2_980(g31297,g30144,g27837);
  AN2 AND2_981(g27183,g26055,g16658);
  AN2 AND2_982(g33376,g32294,g21268);
  AN2 AND2_983(g27673,g25769,g23541);
  AN2 AND2_984(g22004,g5742,g21562);
  AN2 AND2_985(g23008,g1570,g19783);
  AN2 AND2_986(g33889,g33303,g20641);
  AN4 AND4_65(g11123,g5644,g7028,g5630,g9864);
  AN2 AND2_987(g24464,g3480,g23112);
  AN3 AND3_56(I24027,g3029,g3034,g8426);
  AN2 AND2_988(g16885,g6605,g14950);
  AN2 AND2_989(g32169,g31014,g23046);
  AN2 AND2_990(g18575,g2878,g16349);
  AN2 AND2_991(g18474,g2287,g15224);
  AN2 AND2_992(g29902,g28430,g23377);
  AN2 AND2_993(g30289,g28884,g24000);
  AN2 AND2_994(g29377,g28132,g19387);
  AN2 AND2_995(g13807,g4504,g10606);
  AN2 AND2_996(g18711,g15136,g15915);
  AN2 AND2_997(g32168,g30597,g25185);
  AN2 AND2_998(g32410,g4933,g30997);
  AN4 AND4_66(g28991,g14438,g25209,g26424,g27469);
  AN2 AND2_999(g13974,g6243,g12578);
  AN2 AND2_1000(g18327,g1636,g17873);
  AN2 AND2_1001(g24797,g22872,g19960);
  AN2 AND2_1002(g30023,g28508,g20570);
  AN2 AND2_1003(g21712,g294,g20283);
  AN3 AND3_57(I24482,g9364,g9607,g5057);
  AN2 AND2_1004(g18109,g437,g17015);
  AN2 AND2_1005(g27508,g26549,g17684);
  AN2 AND2_1006(g16763,g6239,g14937);
  AN2 AND2_1007(g27634,g26805,g26793);
  AN2 AND2_1008(g34309,g13947,g34147);
  AN2 AND2_1009(g21914,g5077,g21468);
  AN2 AND2_1010(g24292,g4443,g22550);
  AN2 AND2_1011(g30224,g28704,g23896);
  AN2 AND2_1012(g18537,g6856,g15277);
  AN4 AND4_67(I24710,g24071,g24072,g24073,g24074);
  AN2 AND2_1013(g34224,g33736,g22670);
  AN3 AND3_58(g30308,g29178,g7004,g5297);
  AN2 AND2_1014(g22106,g6497,g18833);
  AN3 AND3_59(I24552,g9733,g9316,g5747);
  AN2 AND2_1015(g29645,g1714,g29018);
  AN3 AND3_60(I24003,g8097,g8334,g3045);
  AN4 AND4_68(g17613,g11547,g11592,g11640,I18568);
  AN2 AND2_1016(g34571,g27225,g34299);
  AN2 AND2_1017(g18108,g433,g17015);
  AN2 AND2_1018(g14207,g8639,g11793);
  AN2 AND2_1019(g21907,g5033,g21468);
  AN4 AND4_69(I31286,g30825,g31846,g32868,g32869);
  AN3 AND3_61(I13862,g7232,g7219,g7258);
  AN2 AND2_1020(g15077,g2138,g12955);
  AN2 AND2_1021(g24409,g3484,g23112);
  AN2 AND2_1022(g25966,g9364,g24985);
  AN4 AND4_70(I31306,g30614,g31850,g32896,g32897);
  AN2 AND2_1023(g13265,g9018,g11493);
  AN2 AND2_1024(g18283,g1384,g16136);
  AN2 AND2_1025(g15706,g13296,g13484);
  AN2 AND2_1026(g18606,g3133,g16987);
  AN2 AND2_1027(g18492,g2523,g15426);
  AN2 AND2_1028(g18303,g1536,g16489);
  AN2 AND2_1029(g24408,g23989,g18946);
  AN2 AND2_1030(g24635,g19874,g22883);
  AN2 AND2_1031(g34495,g34274,g19365);
  AN2 AND2_1032(g22033,g5925,g19147);
  AN2 AND2_1033(g27213,g26026,g16721);
  AN2 AND2_1034(g18750,g15145,g17847);
  AN2 AND2_1035(g31520,g29879,g23507);
  AN4 AND4_71(I31187,g32726,g32727,g32728,g32729);
  AN3 AND3_62(g33520,g32888,I31296,I31297);
  AN2 AND2_1036(g18982,g3835,g16159);
  AN2 AND2_1037(g18381,g1882,g15171);
  AN2 AND2_1038(g34687,g14181,g34543);
  AN2 AND2_1039(g21941,g5232,g18997);
  AN2 AND2_1040(g26842,g2894,g24522);
  AN3 AND3_63(I27429,g25562,g26424,g22698);
  AN2 AND2_1041(g27452,g26400,g17600);
  AN2 AND2_1042(g21382,g10086,g17625);
  AN2 AND2_1043(g29632,g28899,g22417);
  AN2 AND2_1044(g31211,g10156,g30102);
  AN4 AND4_72(g26195,g25357,g6856,g11709,g7558);
  AN2 AND2_1045(g34752,g34675,g19544);
  AN2 AND2_1046(g23675,g19050,g9104);
  AN2 AND2_1047(g18174,g739,g17328);
  AN2 AND2_1048(g27311,g12431,g26693);
  AN2 AND2_1049(g18796,g6167,g15348);
  AN2 AND2_1050(g28725,g27596,g20779);
  AN2 AND2_1051(g32084,g10948,g30825);
  AN2 AND2_1052(g32110,g31639,g29921);
  AN2 AND2_1053(g16596,g5941,g14892);
  AN2 AND2_1054(g28114,g25869,g27051);
  AN2 AND2_1055(g25571,I24694,I24695);
  AN2 AND2_1056(g33860,g33270,g20501);
  AN2 AND2_1057(g32321,g27613,g31376);
  AN2 AND2_1058(g16243,g6483,g14275);
  AN2 AND2_1059(g29661,g1687,g29015);
  AN2 AND2_1060(g29547,g1748,g28857);
  AN2 AND2_1061(g29895,g2495,g29170);
  AN2 AND2_1062(g28107,g27970,g18874);
  AN2 AND2_1063(g10683,g7289,g4438);
  AN2 AND2_1064(g32179,g31748,g27907);
  AN2 AND2_1065(g21935,g5196,g18997);
  AN2 AND2_1066(g18390,g1978,g15171);
  AN2 AND2_1067(g31497,g20041,g29930);
  AN3 AND3_64(g33497,g32723,I31181,I31182);
  AN2 AND2_1068(g20109,g17954,g17616);
  AN2 AND2_1069(g24327,g4549,g22228);
  AN2 AND2_1070(g21883,g4141,g19801);
  AN2 AND2_1071(g32178,g31747,g27886);
  AN2 AND2_1072(g15876,g13512,g13223);
  AN2 AND2_1073(g24537,g22626,g10851);
  AN2 AND2_1074(g11116,g9960,g6466);
  AN2 AND2_1075(g20108,g15508,g11048);
  AN2 AND2_1076(g34842,g34762,g20168);
  AN2 AND2_1077(g18192,g817,g17821);
  AN2 AND2_1078(g22012,g5752,g21562);
  AN2 AND2_1079(g26544,g7446,g24357);
  AN4 AND4_73(I27504,g24077,g24078,g24079,g24080);
  AN3 AND3_65(I18620,g13156,g11450,g11498);
  AN2 AND2_1080(g25816,g8164,g24604);
  AN2 AND2_1081(g33700,g33148,g11012);
  AN2 AND2_1082(g33126,g9044,g32201);
  AN2 AND2_1083(g31987,g31767,g22198);
  AN2 AND2_1084(g29551,g2173,g28867);
  AN2 AND2_1085(g29572,g1620,g28885);
  AN2 AND2_1086(g26713,g25447,g20714);
  AN4 AND4_74(I31217,g32768,g32769,g32770,g32771);
  AN2 AND2_1087(g34489,g34421,g19068);
  AN2 AND2_1088(g24283,g4411,g22550);
  AN2 AND2_1089(g18522,g2671,g15509);
  AN2 AND2_1090(g27350,g10217,g26803);
  AN2 AND2_1091(g18663,g4311,g17367);
  AN2 AND2_1092(g24606,g5489,g23630);
  AN2 AND2_1093(g25976,g9443,g25000);
  AN2 AND2_1094(g24303,g4369,g22228);
  AN2 AND2_1095(g16670,g5953,g14999);
  AN2 AND2_1096(g27820,g7670,g25932);
  AN2 AND2_1097(g34525,g34297,g19528);
  AN4 AND4_75(g28141,g10831,g11797,g11261,g27163);
  AN2 AND2_1098(g34488,g34417,g18988);
  AN2 AND2_1099(g28652,g27282,g10288);
  AN2 AND2_1100(g13493,g9880,g11866);
  AN3 AND3_66(g25374,g5366,g23789,I24527);
  AN2 AND2_1101(g31943,g4717,g30614);
  AN3 AND3_67(I24505,g9607,g9229,g5057);
  AN2 AND2_1102(g21729,g3021,g20330);
  AN2 AND2_1103(g26610,g14198,g24405);
  AN2 AND2_1104(g33339,g32221,g20634);
  AN2 AND2_1105(g33943,g33384,g21609);
  AN2 AND2_1106(g31296,g30119,g27779);
  AN2 AND2_1107(g34558,g34353,g20578);
  AN2 AND2_1108(g16734,g5961,g14735);
  AN2 AND2_1109(g23577,g19444,g13033);
  AN2 AND2_1110(g18483,g2453,g15426);
  AN2 AND2_1111(g24750,g17662,g22472);
  AN2 AND2_1112(g32334,g31375,g23568);
  AN2 AND2_1113(g21728,g3010,g20330);
  AN2 AND2_1114(g33338,g32220,g20633);
  AN2 AND2_1115(g28263,g23747,g27711);
  AN2 AND2_1116(g16930,g239,g13132);
  AN2 AND2_1117(g23439,g13771,g20452);
  AN2 AND2_1118(g11035,g5441,g9800);
  AN2 AND2_1119(g18553,g2827,g15277);
  AN2 AND2_1120(g13035,g8497,g11033);
  AN2 AND2_1121(g26270,g1700,g25275);
  AN2 AND2_1122(g31969,g31189,g22139);
  AN2 AND2_1123(g29784,g28331,g23247);
  AN2 AND2_1124(g26124,g1811,g25116);
  AN2 AND2_1125(g22920,g19764,g19719);
  AN2 AND2_1126(g16667,g5268,g14659);
  AN2 AND2_1127(g20174,g5503,g17754);
  AN2 AND2_1128(g29376,g14002,g28504);
  AN2 AND2_1129(g27413,g26576,g17530);
  AN2 AND2_1130(g34865,g16540,g34836);
  AN2 AND2_1131(g16965,g269,g13140);
  AN2 AND2_1132(g18949,g10183,g17625);
  AN2 AND2_1133(g31968,g31757,g22168);
  AN2 AND2_1134(g18326,g1664,g17873);
  AN2 AND2_1135(g24796,g7097,g23714);
  AN2 AND2_1136(g11142,g6381,g10207);
  AN2 AND2_1137(g27691,g25778,g23609);
  AN4 AND4_76(g17724,g11547,g11592,g11640,I18713);
  AN2 AND2_1138(g29354,g4961,g28421);
  AN4 AND4_77(I27533,g21143,g24125,g24126,g24127);
  AN2 AND2_1139(g18536,g2748,g15277);
  AN2 AND2_1140(g23349,g13662,g20182);
  AN2 AND2_1141(g22121,g6593,g19277);
  AN2 AND2_1142(g29888,g28418,g23352);
  AN2 AND2_1143(g33855,g33265,g20441);
  AN2 AND2_1144(g14206,g8655,g11790);
  AN2 AND2_1145(g21906,g5022,g21468);
  AN2 AND2_1146(g18702,g15133,g16856);
  AN2 AND2_1147(g21348,g10121,g17625);
  AN2 AND2_1148(g18757,g5352,g15595);
  AN2 AND2_1149(g31527,g7553,g29343);
  AN2 AND2_1150(g23083,g16076,g19878);
  AN2 AND2_1151(g23348,g15570,g21393);
  AN2 AND2_1152(g15076,g2130,g12955);
  AN2 AND2_1153(g33870,g33280,g20545);
  AN2 AND2_1154(g33411,g32361,g21410);
  AN3 AND3_68(g33527,g32939,I31331,I31332);
  AN2 AND2_1155(g26294,g4245,g25230);
  AN4 AND4_78(I31321,g31376,g31852,g32919,g32920);
  AN2 AND2_1156(g16619,g6629,g14947);
  AN2 AND2_1157(g30042,g29142,g12601);
  AN2 AND2_1158(g18252,g990,g16897);
  AN2 AND2_1159(g18621,g3476,g17062);
  AN2 AND2_1160(g25559,g13004,g22649);
  AN2 AND2_1161(g30255,g28748,g23946);
  AN3 AND3_69(g25488,g6404,g23865,I24603);
  AN4 AND4_79(g28833,g21434,g26424,g25388,g27469);
  AN2 AND2_1162(g16618,g6609,g15039);
  AN2 AND2_1163(g34679,g14093,g34539);
  AN2 AND2_1164(g18564,g2844,g16349);
  AN2 AND2_1165(g30188,g28644,g23841);
  AN2 AND2_1166(g24192,g311,g22722);
  AN2 AND2_1167(g30124,g28580,g21055);
  AN2 AND2_1168(g16279,g4512,g14424);
  AN2 AND2_1169(g34678,g34490,g19431);
  AN2 AND2_1170(g27020,g4601,g25852);
  AN2 AND2_1171(g31503,g20041,g29945);
  AN3 AND3_70(I18716,g13156,g11450,g6756);
  AN4 AND4_80(I31186,g31376,g31828,g32724,g32725);
  AN3 AND3_71(g33503,g32765,I31211,I31212);
  AN2 AND2_1172(g24663,g16621,g22974);
  AN2 AND2_1173(g33867,g33277,g20529);
  AN2 AND2_1174(g17682,g9742,g14637);
  AN2 AND2_1175(g34686,g34494,g19494);
  AN2 AND2_1176(g13523,g7046,g12246);
  AN2 AND2_1177(g18183,g781,g17328);
  AN2 AND2_1178(g18673,g4643,g15758);
  AN2 AND2_1179(g25865,g25545,g18991);
  AN4 AND4_81(g26218,g25357,g6856,g7586,g11686);
  AN2 AND2_1180(g18397,g2004,g15373);
  AN2 AND2_1181(g30030,g29198,g12347);
  AN2 AND2_1182(g30267,g28776,g23967);
  AN3 AND3_72(g34093,g20114,g33755,g9104);
  AN2 AND2_1183(g33450,g32266,g29737);
  AN2 AND2_1184(g22760,g9360,g20237);
  AN2 AND2_1185(g22134,g6653,g19277);
  AN2 AND2_1186(g27113,g25997,g16522);
  AN2 AND2_1187(g32242,g31245,g20324);
  AN2 AND2_1188(g18509,g2587,g15509);
  AN2 AND2_1189(g22029,g5901,g19147);
  AN2 AND2_1190(g31707,g30081,g23886);
  AN2 AND2_1191(g34065,g33813,g23148);
  AN3 AND3_73(g33819,g23088,g33176,g9104);
  AN2 AND2_1192(g33707,g33174,g13346);
  AN2 AND2_1193(g18933,g16237,g13597);
  AN2 AND2_1194(g33910,g33134,g7836);
  AN2 AND2_1195(g24553,g22983,g19539);
  AN2 AND2_1196(g26160,g2453,g25138);
  AN2 AND2_1197(g28273,g27927,g23729);
  AN2 AND2_1198(g7696,g2955,g2950);
  AN2 AND2_1199(g18508,g2606,g15509);
  AN2 AND2_1200(g22028,g5893,g19147);
  AN2 AND2_1201(g27302,g1848,g26680);
  AN2 AND2_1202(g18634,g3813,g17096);
  AN2 AND2_1203(g21333,g1300,g15740);
  AN2 AND2_1204(g23415,g20077,g20320);
  AN2 AND2_1205(g27357,g26400,g17414);
  AN2 AND2_1206(g25042,g23262,g20496);
  AN2 AND2_1207(g31496,g2338,g30312);
  AN2 AND2_1208(g33818,g33236,g20113);
  AN2 AND2_1209(g24949,g23796,g20751);
  AN3 AND3_74(g33496,g32714,I31176,I31177);
  AN2 AND2_1210(g19461,g11708,g16846);
  AN2 AND2_1211(g27105,g26026,g16511);
  AN2 AND2_1212(g24326,g4552,g22228);
  AN2 AND2_1213(g30219,g28698,g23887);
  AN2 AND2_1214(g17134,g5619,g14851);
  AN2 AND2_1215(g21852,g3909,g21070);
  AN2 AND2_1216(g15839,g3929,g13990);
  AN2 AND2_1217(g34875,g34836,g20073);
  AN2 AND2_1218(g28812,g26972,g13037);
  AN2 AND2_1219(g33111,g24005,g32421);
  AN2 AND2_1220(g34219,g33736,g22942);
  AN2 AND2_1221(g31070,g29814,g25985);
  AN2 AND2_1222(g19145,g8450,g16200);
  AN2 AND2_1223(g24536,g19516,g22635);
  AN2 AND2_1224(g29860,g28389,g23312);
  AN2 AND2_1225(g17506,g9744,g14505);
  AN2 AND2_1226(g25124,g4917,g22908);
  AN2 AND2_1227(g15694,g457,g13437);
  AN2 AND2_1228(g15838,g3602,g14133);
  AN2 AND2_1229(g21963,g5436,g21514);
  AN2 AND2_1230(g24702,g17464,g22342);
  AN2 AND2_1231(g34218,g33744,g22670);
  AN2 AND2_1232(g24757,g7004,g23563);
  AN2 AND2_1233(g31986,g31766,g22197);
  AN2 AND2_1234(g19736,g12136,g17136);
  AN2 AND2_1235(g24904,g11761,g23279);
  AN2 AND2_1236(g28234,g27877,g26686);
  AN2 AND2_1237(g32293,g2827,g30593);
  AN4 AND4_82(I31216,g30937,g31834,g32766,g32767);
  AN2 AND2_1238(g25939,g24583,g19490);
  AN2 AND2_1239(g26277,g2547,g25400);
  AN2 AND2_1240(g18213,g952,g15979);
  AN2 AND2_1241(g32265,g2799,g30567);
  AN2 AND2_1242(g25030,g23251,g20432);
  AN2 AND2_1243(g25938,g8997,g24953);
  AN2 AND2_1244(g25093,g12831,g23493);
  AN2 AND2_1245(g31067,g29484,g22868);
  AN2 AND2_1246(g24564,g23198,g21163);
  AN2 AND2_1247(g29625,g28514,g14226);
  AN3 AND3_75(g29987,g29197,g26424,g22763);
  AN2 AND2_1248(g19393,g691,g16325);
  AN2 AND2_1249(g16884,g6159,g14321);
  AN2 AND2_1250(g18574,g2882,g16349);
  AN2 AND2_1251(g23484,g20160,g20541);
  AN2 AND2_1252(g18452,g2311,g15224);
  AN2 AND2_1253(g18205,g904,g15938);
  AN2 AND2_1254(g31150,g1682,g30063);
  AN2 AND2_1255(g23554,g20390,g13024);
  AN4 AND4_83(I31117,g32624,g32625,g32626,g32627);
  AN2 AND2_1256(g18311,g1554,g16931);
  AN2 AND2_1257(g33801,g33437,g25327);
  AN2 AND2_1258(g24673,g22659,g19748);
  AN2 AND2_1259(g33735,g33118,g19553);
  AN2 AND2_1260(g33877,g33287,g20563);
  AN3 AND3_76(I24582,g9809,g9397,g6093);
  AN2 AND2_1261(g30915,g29886,g24778);
  AN2 AND2_1262(g29943,g2165,g28765);
  AN2 AND2_1263(g34470,g7834,g34325);
  AN2 AND2_1264(g16666,g5200,g14794);
  AN2 AND2_1265(g25875,g8390,g24809);
  AN2 AND2_1266(g31019,g29481,g22856);
  AN3 AND3_77(I18765,g13156,g11450,g11498);
  AN2 AND2_1267(g29644,g28216,g19794);
  AN2 AND2_1268(g29338,g29145,g22181);
  AN2 AND2_1269(g30277,g28817,g23987);
  AN2 AND2_1270(g13063,g8567,g10808);
  AN2 AND2_1271(g31018,g29480,g22855);
  AN2 AND2_1272(g32014,g8715,g30673);
  AN2 AND2_1273(g29969,g28121,g20509);
  AN2 AND2_1274(g30075,g28525,g20662);
  AN2 AND2_1275(g26155,g1945,g25134);
  AN2 AND2_1276(g14221,g8686,g11823);
  AN2 AND2_1277(g21921,g5109,g21468);
  AN2 AND2_1278(g26822,g24841,g13116);
  AN4 AND4_84(I31242,g32805,g32806,g32807,g32808);
  AN4 AND4_85(g16486,g6772,g11592,g6789,I17692);
  AN2 AND2_1279(g18592,g2994,g16349);
  AN2 AND2_1280(g23921,g19379,g4146);
  AN2 AND2_1281(g18756,g5348,g15595);
  AN2 AND2_1282(g34075,g33692,g19517);
  AN2 AND2_1283(g31526,g22521,g29342);
  AN2 AND2_1284(g24634,g22634,g19685);
  AN2 AND2_1285(g30595,g18911,g29847);
  AN3 AND3_78(g33526,g32932,I31326,I31327);
  AN2 AND2_1286(g24872,g23088,g9104);
  AN2 AND2_1287(g29968,g2433,g28843);
  AN2 AND2_1288(g21745,g3017,g20330);
  AN2 AND2_1289(g18780,g5827,g18065);
  AN2 AND2_1290(g12027,g9499,g9729);
  AN2 AND2_1291(g14613,g10602,g10585);
  AN2 AND2_1292(g27249,g25929,g19678);
  AN2 AND2_1293(g21799,g3530,g20924);
  AN2 AND2_1294(g29855,g2287,g29093);
  AN2 AND2_1295(g17770,g7863,g13189);
  AN2 AND2_1296(g21813,g3590,g20924);
  AN2 AND2_1297(g23799,g14911,g21279);
  AN2 AND2_1298(g27482,g26488,g17641);
  AN2 AND2_1299(g15815,g3594,g14075);
  AN2 AND2_1300(g28541,g27403,g20274);
  AN2 AND2_1301(g10947,g9200,g1430);
  AN2 AND2_1302(g18350,g1779,g17955);
  AN3 AND3_79(I24603,g9892,g9467,g6439);
  AN2 AND2_1303(g33402,g32351,g21395);
  AN2 AND2_1304(g29870,g2421,g29130);
  AN2 AND2_1305(g29527,g28945,g22432);
  AN2 AND2_1306(g27710,g26422,g20904);
  AN2 AND2_1307(g21798,g3522,g20924);
  AN2 AND2_1308(g34782,g34711,g33888);
  AN4 AND4_86(I27529,g28038,g24121,g24122,g24123);
  AN2 AND2_1309(g18820,g15166,g15563);
  AN2 AND2_1310(g26853,g94,g24533);
  AN4 AND4_87(g28789,g21434,g26424,g25340,g27440);
  AN2 AND2_1311(g21973,g5511,g19074);
  AN2 AND2_1312(g32116,g31658,g29929);
  AN2 AND2_1313(g27204,g26026,g16689);
  AN2 AND2_1314(g33866,g33276,g20528);
  AN2 AND2_1315(g22899,g19486,g19695);
  AN2 AND2_1316(g21805,g3550,g20924);
  AN2 AND2_1317(g22990,g19555,g19760);
  AN4 AND4_88(I27528,g20998,g24118,g24119,g24120);
  AN2 AND2_1318(g18152,g613,g17533);
  AN2 AND2_1319(g25915,g24926,g9602);
  AN2 AND2_1320(g32041,g13913,g31262);
  AN2 AND2_1321(g18396,g2008,g15373);
  AN2 AND2_1322(g22633,g19359,g19479);
  AN4 AND4_89(g17767,g6772,g11592,g6789,I18765);
  AN2 AND2_1323(g18731,g15140,g16861);
  AN2 AND2_1324(g30266,g28775,g23966);
  AN2 AND2_1325(g28535,g11981,g27088);
  AN2 AND2_1326(g15937,g11950,g14387);
  AN2 AND2_1327(g25201,g12346,g23665);
  AN2 AND2_1328(g22191,g8119,g19875);
  AN2 AND2_1329(g16179,g6187,g14321);
  AN2 AND2_1330(g29867,g1996,g29117);
  AN2 AND2_1331(g29894,g2070,g29169);
  AN2 AND2_1332(g19069,g8397,g16186);
  AN2 AND2_1333(g21732,g3004,g20330);
  AN2 AND2_1334(g16531,g5232,g14656);
  AN2 AND2_1335(g13542,g10053,g11927);
  AN2 AND2_1336(g21934,g5220,g18997);
  AN2 AND2_1337(g18413,g2089,g15373);
  AN2 AND2_1338(g24912,g23687,g20682);
  AN2 AND2_1339(g26119,g11944,g25109);
  AN2 AND2_1340(g24311,g4498,g22228);
  AN2 AND2_1341(g16178,g5845,g14297);
  AN2 AND2_1342(g18691,g4727,g16053);
  AN2 AND2_1343(g15884,g3901,g14113);
  AN2 AND2_1344(g33689,g33144,g11006);
  AN2 AND2_1345(g32340,g31468,g23585);
  AN2 AND2_1346(g29581,g28462,g11796);
  AN2 AND2_1347(g32035,g4176,g30937);
  AN2 AND2_1348(g31280,g29717,g23305);
  AN2 AND2_1349(g17191,g1384,g13242);
  AN2 AND2_1350(g17719,g9818,g14675);
  AN2 AND2_1351(g21761,g3215,g20785);
  AN3 AND3_80(g29315,g29188,g7051,g5990);
  AN4 AND4_90(g27999,g23032,g26200,g26424,g25529);
  AN2 AND2_1352(g26864,g2907,g24548);
  AN2 AND2_1353(g26022,g25271,g20751);
  AN2 AND2_1354(g13436,g9721,g11811);
  AN2 AND2_1355(g18405,g2040,g15373);
  AN2 AND2_1356(g31300,g30148,g27858);
  AN2 AND2_1357(g30167,g28622,g23793);
  AN2 AND2_1358(g30194,g28651,g23849);
  AN2 AND2_1359(g30589,g18898,g29811);
  AN4 AND4_91(I24690,g24043,g24044,g24045,g24046);
  AN3 AND3_81(I24549,g5385,g5390,g9792);
  AN2 AND2_1360(g26749,g24494,g23578);
  AN2 AND2_1361(g27090,g25997,g16423);
  AN3 AND3_82(g29202,g24088,I27508,I27509);
  AN2 AND2_1362(g25782,g2936,g24571);
  AN2 AND2_1363(g32142,g31616,g29965);
  AN2 AND2_1364(g13320,g417,g11048);
  AN2 AND2_1365(g26313,g12645,g25326);
  AN3 AND3_83(g28291,g7411,g2070,g27469);
  AN2 AND2_1366(g29979,g23655,g28991);
  AN2 AND2_1367(g34588,g26082,g34323);
  AN2 AND2_1368(g22861,g19792,g19670);
  AN2 AND2_1369(g27651,g22448,g25781);
  AN2 AND2_1370(g34524,g9083,g34359);
  AN2 AND2_1371(g33102,g32399,g18978);
  AN4 AND4_92(I31007,g32466,g32467,g32468,g32469);
  AN2 AND2_1372(g26276,g2461,g25476);
  AN2 AND2_1373(g26285,g1834,g25300);
  AN2 AND2_1374(g34401,g34199,g21383);
  AN2 AND2_1375(g34477,g26344,g34328);
  AN2 AND2_1376(g22045,g6069,g21611);
  AN2 AND2_1377(g18583,g2936,g16349);
  AN2 AND2_1378(g29590,g2625,g28615);
  AN3 AND3_84(g34119,g20516,g9104,g33755);
  AN2 AND2_1379(g26254,g2413,g25349);
  AN2 AND2_1380(g31066,g29483,g22865);
  AN2 AND2_1381(g31231,g30290,g25239);
  AN2 AND2_1382(g29986,g28468,g23473);
  AN2 AND2_1383(g22099,g6462,g18833);
  AN2 AND2_1384(g27932,g25944,g19369);
  AN2 AND2_1385(g27331,g10177,g26754);
  AN2 AND2_1386(g30118,g28574,g21050);
  AN2 AND2_1387(g24820,g13944,g23978);
  AN2 AND2_1388(g26808,g25521,g21185);
  AN2 AND2_1389(g16762,g5901,g14930);
  AN2 AND2_1390(g20152,g11545,g16727);
  AN2 AND2_1391(g22534,g8766,g21389);
  AN3 AND3_85(g29384,g26424,g22763,g28179);
  AN2 AND2_1392(g22098,g6459,g18833);
  AN2 AND2_1393(g32193,g30732,g25410);
  AN4 AND4_93(I31116,g31154,g31816,g32622,g32623);
  AN3 AND3_86(g24846,g3361,g23555,I24018);
  AN2 AND2_1394(g26101,g1760,g25098);
  AN2 AND2_1395(g33876,g33286,g20562);
  AN2 AND2_1396(g33885,g33296,g20609);
  AN2 AND2_1397(g26177,g2079,g25154);
  AN2 AND2_1398(g18113,g405,g17015);
  AN2 AND2_1399(g18787,g15158,g15634);
  AN2 AND2_1400(g32165,g31669,g27742);
  AN2 AND2_1401(g24731,g6519,g23733);
  AN4 AND4_94(I31041,g31566,g31803,g32513,g32514);
  AN2 AND2_1402(g18282,g1379,g16136);
  AN2 AND2_1403(g34748,g34672,g19529);
  AN2 AND2_1404(g27505,g26519,g17681);
  AN2 AND2_1405(g27404,g26400,g17518);
  AN2 AND2_1406(g31763,g30127,g23965);
  AN2 AND2_1407(g18302,g1514,g16489);
  AN3 AND3_87(g33511,g32823,I31251,I31252);
  AN2 AND2_1408(g15084,g2710,g12983);
  AN2 AND2_1409(g18357,g1816,g17955);
  AN2 AND2_1410(g19545,g3147,g16769);
  AN2 AND2_1411(g29877,g28405,g23340);
  AN2 AND2_1412(g15110,g4245,g14454);
  AN2 AND2_1413(g18105,g417,g17015);
  AN2 AND2_1414(g10724,g3689,g8728);
  AN2 AND2_1415(g22032,g5921,g19147);
  AN2 AND2_1416(g30254,g28747,g23944);
  AN2 AND2_1417(g18743,g5115,g17847);
  AN2 AND2_1418(g27212,g25997,g16717);
  AN2 AND2_1419(g10829,g7289,g4375);
  AN4 AND4_95(I31237,g32798,g32799,g32800,g32801);
  AN2 AND2_1420(g21771,g3255,g20785);
  AN2 AND2_1421(g10828,g6888,g7640);
  AN2 AND2_1422(g18640,g3835,g17096);
  AN2 AND2_1423(g18769,g15151,g18062);
  AN2 AND2_1424(g22061,g6065,g21611);
  AN2 AND2_1425(g30101,g28551,g20780);
  AN2 AND2_1426(g30177,g28631,g23814);
  AN2 AND2_1427(g29526,g28938,g22384);
  AN2 AND2_1428(g17140,g8616,g12968);
  AN2 AND2_1429(g26630,g7592,g24419);
  AN2 AND2_1430(g34560,g34366,g17366);
  AN2 AND2_1431(g18768,g5503,g17929);
  AN2 AND2_1432(g18803,g15161,g15480);
  AN2 AND2_1433(g31480,g1644,g30296);
  AN4 AND4_96(I31142,g32661,g32662,g32663,g32664);
  AN3 AND3_88(g33480,g32600,I31096,I31097);
  AN2 AND2_1434(g24929,g23751,g20875);
  AN2 AND2_1435(g22871,g9523,g20871);
  AN4 AND4_97(g26166,g25357,g11724,g11709,g7558);
  AN2 AND2_1436(g27723,g26512,g21049);
  AN2 AND2_1437(g15654,g3845,g13584);
  AN2 AND2_1438(g31314,g30183,g27937);
  AN2 AND2_1439(g28240,g27356,g17239);
  AN2 AND2_1440(g27149,g25997,g16623);
  AN2 AND2_1441(g30064,g28517,g20630);
  AN4 AND4_98(g17766,g6772,g11592,g11640,I18762);
  AN2 AND2_1442(g27433,g26519,g17583);
  AN2 AND2_1443(g27387,g26488,g17499);
  AN2 AND2_1444(g15936,g475,g13999);
  AN2 AND2_1445(g25285,g22152,g13061);
  AN2 AND2_1446(g29866,g1906,g29116);
  AN2 AND2_1447(g27148,g25997,g16622);
  AN2 AND2_1448(g21882,g4057,g19801);
  AN2 AND2_1449(g21991,g5595,g19074);
  AN2 AND2_1450(g26485,g24968,g10502);
  AN2 AND2_1451(g23991,g19209,g21428);
  AN2 AND2_1452(g27097,g25867,g22526);
  AN2 AND2_1453(g33721,g33163,g19440);
  AN2 AND2_1454(g19656,g2807,g15844);
  AN2 AND2_1455(g27104,g25997,g16510);
  AN2 AND2_1456(g16751,g13155,g13065);
  AN2 AND2_1457(g16807,g6585,g14978);
  AN2 AND2_1458(g27646,g13094,g25773);
  AN2 AND2_1459(g25900,g24390,g19368);
  AN2 AND2_1460(g34874,g34833,g20060);
  AN2 AND2_1461(g23407,g9295,g20273);
  AN2 AND2_1462(g33243,g32124,g19947);
  AN2 AND2_1463(g28563,g11981,g27100);
  AN2 AND2_1464(g25466,g23574,g21346);
  AN2 AND2_1465(g19680,g12028,g17013);
  AN2 AND2_1466(g33431,g32364,g32377);
  AN2 AND2_1467(g16639,g6291,g14974);
  AN2 AND2_1468(g26712,g24508,g24463);
  AN3 AND3_89(I17741,g14988,g11450,g11498);
  AN2 AND2_1469(g18662,g15126,g17367);
  AN2 AND2_1470(g32175,g31709,g27858);
  AN2 AND2_1471(g30166,g28621,g23792);
  AN2 AND2_1472(g30009,g29034,g10518);
  AN2 AND2_1473(g24302,g15124,g22228);
  AN2 AND2_1474(g16638,g6271,g14773);
  AN2 AND2_1475(g33269,g31970,g15582);
  AN2 AND2_1476(g34665,g34583,g19067);
  AN3 AND3_90(g22472,g7753,g9285,g21289);
  AN2 AND2_1477(g18890,g10158,g17625);
  AN2 AND2_1478(g13492,g9856,g11865);
  AN2 AND2_1479(g27369,g25894,g25324);
  AN2 AND2_1480(g24743,g22708,g19789);
  AN2 AND2_1481(g30008,g29191,g12297);
  AN2 AND2_1482(g18249,g1216,g16897);
  AN2 AND2_1483(g33942,g33383,g21608);
  AN2 AND2_1484(g33341,g32223,g20640);
  AN2 AND2_1485(g18482,g2472,g15426);
  AN2 AND2_1486(g14506,g1430,g10755);
  AN2 AND2_1487(g29688,g2509,g28713);
  AN4 AND4_99(I31006,g31376,g31796,g32464,g32465);
  AN2 AND2_1488(g29624,g28491,g8070);
  AN2 AND2_1489(g14028,g8673,g11797);
  AN2 AND2_1490(g18248,g15067,g16897);
  AN2 AND2_1491(g16841,g5913,g14858);
  AN2 AND2_1492(g18710,g15135,g17302);
  AN2 AND2_1493(g34476,g34399,g18891);
  AN2 AND2_1494(g34485,g34411,g18952);
  AN2 AND2_1495(g18552,g2815,g15277);
  AN2 AND2_1496(g24640,g6509,g23733);
  AN2 AND2_1497(g24769,g19619,g23058);
  AN2 AND2_1498(g19631,g1484,g16093);
  AN2 AND2_1499(g18204,g914,g15938);
  AN4 AND4_100(I31222,g32775,g32776,g32777,g32778);
  AN2 AND2_1500(g27412,g26576,g17529);
  AN2 AND2_1501(g34555,g34349,g20512);
  AN2 AND2_1502(g18779,g5821,g18065);
  AN2 AND2_1503(g22071,g6251,g19210);
  AN2 AND2_1504(g24803,g22901,g20005);
  AN3 AND3_91(g33734,g7806,g33136,I31593);
  AN2 AND2_1505(g30914,g29873,g20887);
  AN2 AND2_1506(g21759,g3199,g20785);
  AN2 AND2_1507(g15117,g4300,g14454);
  AN2 AND2_1508(g23725,g14772,g21138);
  AN2 AND2_1509(g18778,g5817,g18065);
  AN2 AND2_1510(g25874,g11118,g24665);
  AN2 AND2_1511(g27229,g26055,g16774);
  AN2 AND2_1512(g31993,g31774,g22214);
  AN2 AND2_1513(g21758,g3191,g20785);
  AN2 AND2_1514(g26176,g1964,g25467);
  AN2 AND2_1515(g26092,g9766,g25083);
  AN2 AND2_1516(g18786,g15156,g15345);
  AN2 AND2_1517(g27228,g26055,g16773);
  AN3 AND3_92(g24881,g3050,g23211,I24048);
  AN4 AND4_101(I31347,g32956,g32957,g32958,g32959);
  AN2 AND2_1518(g22859,g9456,g20734);
  AN2 AND2_1519(g26154,g1830,g25426);
  AN2 AND2_1520(g30239,g28728,g23923);
  AN2 AND2_1521(g17785,g13341,g10762);
  AN2 AND2_1522(g25166,g17506,g23571);
  AN2 AND2_1523(g31131,g2393,g30020);
  AN2 AND2_1524(g18647,g4040,g17271);
  AN2 AND2_1525(g34074,g33685,g19498);
  AN2 AND2_1526(g30594,g18898,g29846);
  AN2 AND2_1527(g18356,g1802,g17955);
  AN2 AND2_1528(g29876,g28404,g23339);
  AN2 AND2_1529(g29885,g28416,g23350);
  AN2 AND2_1530(g21744,g3103,g20330);
  AN2 AND2_1531(g30238,g28727,g23922);
  AN2 AND2_1532(g34567,g34377,g17491);
  AN3 AND3_93(I31600,g31009,g8400,g7809);
  AN2 AND2_1533(g28440,g27274,g20059);
  AN2 AND2_1534(g18826,g7097,g15680);
  AN2 AND2_1535(g18380,g1926,g15171);
  AN2 AND2_1536(g19571,g3498,g16812);
  AN3 AND3_94(g33487,g32649,I31131,I31132);
  AN2 AND2_1537(g22172,g8064,g19857);
  AN2 AND2_1538(g29854,g2197,g29092);
  AN2 AND2_1539(g21849,g3889,g21070);
  AN2 AND2_1540(g21940,g5228,g18997);
  AN4 AND4_102(I31236,g30735,g31837,g32796,g32797);
  AN2 AND2_1541(g15814,g3574,g13920);
  AN2 AND2_1542(g31502,g2472,g29311);
  AN2 AND2_1543(g28573,g7349,g27059);
  AN3 AND3_95(g25485,g6098,g22220,I24600);
  AN3 AND3_96(g33502,g32758,I31206,I31207);
  AN2 AND2_1544(g29511,g1736,g28783);
  AN2 AND2_1545(g31210,g2509,g30100);
  AN4 AND4_103(I31351,g30937,g31858,g32961,g32962);
  AN2 AND2_1546(g18233,g1094,g16326);
  AN2 AND2_1547(g28247,g27147,g19675);
  AN2 AND2_1548(g21848,g3913,g21070);
  AN2 AND2_1549(g15807,g3570,g13898);
  AN2 AND2_1550(g18182,g776,g17328);
  AN2 AND2_1551(g27310,g26574,g23059);
  AN2 AND2_1552(g18651,g15102,g16249);
  AN2 AND2_1553(g18672,g15127,g15758);
  AN2 AND2_1554(g34382,g34167,g20618);
  AN2 AND2_1555(g30185,g28640,g23838);
  AN2 AND2_1556(g34519,g34293,g19504);
  AN2 AND2_1557(g17151,g8659,g12996);
  AN2 AND2_1558(g21804,g3542,g20924);
  AN2 AND2_1559(g34185,g33702,g24389);
  AN2 AND2_1560(g27627,g13266,g25790);
  AN2 AND2_1561(g25570,I24689,I24690);
  AN2 AND2_1562(g27959,g25948,g19374);
  AN2 AND2_1563(g28612,g27524,g20539);
  AN3 AND3_97(g34092,g33750,g9104,g18957);
  AN2 AND2_1564(g30154,g28611,g23769);
  AN2 AND2_1565(g28324,g9875,g27687);
  AN2 AND2_1566(g24482,g6875,g23055);
  AN2 AND2_1567(g31278,g29716,g23302);
  AN2 AND2_1568(g34518,g34292,g19503);
  AN2 AND2_1569(g32274,g31256,g20447);
  AN2 AND2_1570(g27050,g25789,g22338);
  AN2 AND2_1571(g27958,g25950,g22449);
  AN2 AND2_1572(g25907,g24799,g22519);
  AN2 AND2_1573(g24710,g22679,g19771);
  AN2 AND2_1574(g27378,g26089,g20052);
  AN4 AND4_104(I31137,g32654,g32655,g32656,g32657);
  AN2 AND2_1575(g18331,g1682,g17873);
  AN3 AND3_98(I27364,g25541,g26424,g22698);
  AN2 AND2_1576(g24552,g22487,g19538);
  AN3 AND3_99(g33469,g32519,I31041,I31042);
  AN2 AND2_1577(g28251,g27826,g23662);
  AN2 AND2_1578(g30935,g8808,g29745);
  AN2 AND2_1579(g28272,g27721,g26548);
  AN2 AND2_1580(g31286,g30159,g27858);
  AN2 AND2_1581(g32122,g31646,g29944);
  AN2 AND2_1582(g18513,g2575,g15509);
  AN2 AND2_1583(g21332,g996,g15739);
  AN2 AND2_1584(g18449,g12852,g15224);
  AN3 AND3_100(I26972,g25011,g26424,g22698);
  AN2 AND2_1585(g27386,g26488,g17498);
  AN2 AND2_1586(g19752,g2771,g15864);
  AN3 AND3_101(g33468,g32512,I31036,I31037);
  AN2 AND2_1587(g15841,g4273,g13868);
  AN2 AND2_1588(g25567,I24674,I24675);
  AN2 AND2_1589(g27096,g26026,g16475);
  AN2 AND2_1590(g18448,g2153,g18008);
  AN2 AND2_1591(g29550,g28990,g22457);
  AN2 AND2_1592(g32034,g14124,g31239);
  AN2 AND2_1593(g25238,g12466,g23732);
  AN2 AND2_1594(g16806,g6247,g14971);
  AN2 AND2_1595(g29314,g29005,g22144);
  AN2 AND2_1596(g22059,g6148,g21611);
  AN2 AND2_1597(g21962,g5428,g21514);
  AN2 AND2_1598(g18505,g2583,g15509);
  AN2 AND2_1599(g21361,g7869,g16066);
  AN2 AND2_1600(g22025,g5905,g19147);
  AN2 AND2_1601(g18404,g2066,g15373);
  AN2 AND2_1602(g24786,g661,g23654);
  AN2 AND2_1603(g33815,g33449,g12911);
  AN2 AND2_1604(g32292,g31269,g20530);
  AN2 AND2_1605(g10898,g3706,g9100);
  AN2 AND2_1606(g18717,g4849,g15915);
  AN2 AND2_1607(g22058,g6098,g21611);
  AN2 AND2_1608(g31187,g10118,g30090);
  AN2 AND2_1609(g32153,g31646,g29999);
  AN2 AND2_1610(g24647,g19903,g22907);
  AN2 AND2_1611(g33677,g33443,g31937);
  AN2 AND2_1612(g31975,g31761,g22177);
  AN4 AND4_105(g13252,g11561,g11511,g11469,g699);
  AN2 AND2_1613(g18212,g947,g15979);
  AN2 AND2_1614(g29596,g27823,g28620);
  AN2 AND2_1615(g24945,g23183,g20197);
  AN3 AND3_102(g10719,g6841,g2138,g2130);
  AN2 AND2_1616(g16517,g5248,g14797);
  AN2 AND2_1617(g21833,g15096,g20453);
  AN2 AND2_1618(g30215,g28690,g23881);
  AN2 AND2_1619(g32409,g4754,g30996);
  AN2 AND2_1620(g14719,g4392,g10830);
  AN2 AND2_1621(g34215,g33778,g22670);
  AN2 AND2_1622(g30577,g26267,g29679);
  AN2 AND2_1623(g34577,g24577,g34307);
  AN3 AND3_103(g25518,g6444,g23865,I24625);
  AN2 AND2_1624(g27428,g26400,g17576);
  AN2 AND2_1625(g13564,g4480,g12820);
  AN2 AND2_1626(g22044,g6058,g21611);
  AN2 AND2_1627(g26304,g2697,g25246);
  AN2 AND2_1628(g31143,g29506,g22999);
  AN4 AND4_106(I24709,g21256,g24068,g24069,g24070);
  AN4 AND4_107(I31021,g31070,g31799,g32485,g32486);
  AN2 AND2_1629(g24998,g17412,g23408);
  AN2 AND2_1630(g12730,g9024,g4349);
  AN2 AND2_1631(g27765,g4146,g25886);
  AN2 AND2_1632(g24651,g2741,g23472);
  AN2 AND2_1633(g24672,g19534,g22981);
  AN2 AND2_1634(g14832,g1489,g10939);
  AN2 AND2_1635(g29773,g28203,g10233);
  AN2 AND2_1636(g27690,g25784,g23607);
  AN2 AND2_1637(g16193,g6533,g14348);
  AN2 AND2_1638(g27549,g26576,g14785);
  AN2 AND2_1639(g31169,g10083,g30079);
  AN2 AND2_1640(g11397,g5360,g7139);
  AN2 AND2_1641(g18723,g4922,g16077);
  AN2 AND2_1642(g25883,g13728,g24699);
  AN2 AND2_1643(g28360,g27401,g19861);
  AN2 AND2_1644(g22120,g6585,g19277);
  AN2 AND2_1645(g33884,g33295,g20590);
  AN2 AND2_1646(g15116,g4297,g14454);
  AN2 AND2_1647(g18149,g608,g17533);
  AN2 AND2_1648(g27548,g26576,g17763);
  AN2 AND2_1649(g31168,g2241,g30077);
  AN2 AND2_1650(g32164,g30733,g25171);
  AN2 AND2_1651(g18433,g2197,g18008);
  AN2 AND2_1652(g33410,g32360,g21409);
  AN2 AND2_1653(g18387,g1955,g15171);
  AN2 AND2_1654(g24331,g6977,g22228);
  AN2 AND2_1655(g30083,g28533,g20698);
  AN2 AND2_1656(g13509,g9951,g11889);
  AN2 AND2_1657(g27504,g26519,g17680);
  AN2 AND2_1658(g18620,g3470,g17062);
  AN2 AND2_1659(g18148,g562,g17533);
  AN2 AND2_1660(g21947,g5256,g18997);
  AN2 AND2_1661(g30284,g28852,g23994);
  AN2 AND2_1662(g34083,g33714,g19573);
  AN2 AND2_1663(g34348,g34125,g20128);
  AN3 AND3_104(I31593,g31003,g8350,g7788);
  AN3 AND3_105(g33479,g32593,I31091,I31092);
  AN2 AND2_1664(g34284,g34046,g19351);
  AN2 AND2_1665(g21605,g13005,g15695);
  AN4 AND4_108(I31346,g31021,g31857,g32954,g32955);
  AN2 AND2_1666(g33363,g32262,g20918);
  AN2 AND2_1667(g13508,g9927,g11888);
  AN2 AND2_1668(g18104,g392,g17015);
  AN2 AND2_1669(g18811,g6500,g15483);
  AN2 AND2_1670(g18646,g4031,g17271);
  AN4 AND4_109(I31122,g32631,g32632,g32633,g32634);
  AN2 AND2_1671(g14612,g11971,g11993);
  AN2 AND2_1672(g31478,g29764,g23410);
  AN2 AND2_1673(g8234,g4515,g4521);
  AN2 AND2_1674(g31015,g29476,g22758);
  AN2 AND2_1675(g18343,g12847,g17955);
  AN3 AND3_106(g24897,g3401,g23223,I24064);
  AN2 AND2_1676(g29839,g1728,g29045);
  AN2 AND2_1677(g30566,g26247,g29507);
  AN3 AND3_107(g33478,g32584,I31086,I31087);
  AN2 AND2_1678(g24961,g23193,g20209);
  AN2 AND2_1679(g21812,g3586,g20924);
  AN2 AND2_1680(g17146,g5965,g14895);
  AN2 AND2_1681(g34566,g34376,g17489);
  AN2 AND2_1682(g28451,g27283,g20090);
  AN2 AND2_1683(g16222,g6513,g14348);
  AN2 AND2_1684(g31486,g29777,g23422);
  AN2 AND2_1685(g32327,g31319,g23544);
  AN2 AND2_1686(g29667,g2671,g29157);
  AN2 AND2_1687(g29838,g1636,g29044);
  AN2 AND2_1688(g27129,g26026,g16584);
  AN3 AND3_108(g33486,g32642,I31126,I31127);
  AN2 AND2_1689(g32109,g31609,g29920);
  AN2 AND2_1690(g21951,g5272,g18997);
  AN2 AND2_1691(g26852,g24975,g24958);
  AN2 AND2_1692(g21972,g15152,g19074);
  AN4 AND4_110(g27057,g7791,g6219,g6227,g26261);
  AN2 AND2_1693(g19610,g1141,g16069);
  AN2 AND2_1694(g18369,g12848,g15171);
  AN2 AND2_1695(g24717,g22684,g19777);
  AN2 AND2_1696(g27128,g25997,g16583);
  AN2 AND2_1697(g28246,g8572,g27976);
  AN4 AND4_111(I31292,g32877,g32878,g32879,g32880);
  AN2 AND2_1698(g32108,g31631,g29913);
  AN2 AND2_1699(g30139,g28596,g21184);
  AN2 AND2_1700(g18368,g1728,g17955);
  AN2 AND2_1701(g34139,g33827,g23314);
  AN2 AND2_1702(g16703,g5889,g15002);
  AN2 AND2_1703(g22632,g19356,g19476);
  AN2 AND2_1704(g31223,g20028,g29689);
  AN2 AND2_1705(g21795,g3506,g20924);
  AN2 AND2_1706(g32283,g31259,g20506);
  AN2 AND2_1707(g27323,g26268,g23086);
  AN2 AND2_1708(g30138,g28595,g21182);
  AN2 AND2_1709(g27299,g26546,g23028);
  AN2 AND2_1710(g29619,g2269,g29060);
  AN2 AND2_1711(g32303,g27550,g31376);
  AN2 AND2_1712(g34138,g33929,g23828);
  AN2 AND2_1713(g11047,g6474,g9212);
  AN2 AND2_1714(g18412,g2098,g15373);
  AN4 AND4_112(I31136,g29385,g32651,g32652,g32653);
  AN2 AND2_1715(g11205,g8217,g8439);
  AN2 AND2_1716(g13047,g8534,g11042);
  AN2 AND2_1717(g27298,g26573,g23026);
  AN2 AND2_1718(g29618,g28870,g22384);
  AN2 AND2_1719(g19383,g16893,g13223);
  AN2 AND2_1720(g34415,g34207,g21458);
  AN2 AND2_1721(g18133,g15055,g17249);
  AN2 AND2_1722(g23514,g20149,g11829);
  AN2 AND2_1723(g26484,g24946,g8841);
  AN2 AND2_1724(g33110,g32404,g32415);
  AN2 AND2_1725(g13912,g5551,g12450);
  AN2 AND2_1726(g34333,g9984,g34192);
  AN2 AND2_1727(g24723,g17490,g22384);
  AN2 AND2_1728(g31321,g30146,g27886);
  AN2 AND2_1729(g18229,g1099,g16326);
  AN2 AND2_1730(g33922,g33448,g7202);
  AN2 AND2_1731(g14061,g8715,g11834);
  AN3 AND3_109(g33531,g32967,I31351,I31352);
  AN2 AND2_1732(g18228,g1061,g16129);
  AN2 AND2_1733(g24387,g3457,g22761);
  AN2 AND2_1734(g26312,g2704,g25264);
  AN2 AND2_1735(g34963,g34946,g23041);
  AN4 AND4_113(g26200,g24688,g10678,g10658,g10627);
  AN2 AND2_1736(g32174,g31708,g27837);
  AN2 AND2_1737(g21163,g16321,g4878);
  AN2 AND2_1738(g21012,g16304,g4688);
  AN2 AND2_1739(g28151,g8426,g27295);
  AN2 AND2_1740(g18716,g4878,g15915);
  AN2 AND2_1741(g31186,g2375,g30088);
  AN2 AND2_1742(g33186,g32037,g22830);
  AN2 AND2_1743(g24646,g22640,g19711);
  AN2 AND2_1744(g33676,g33125,g7970);
  AN2 AND2_1745(g33373,g32288,g21205);
  AN2 AND2_1746(g16516,g5228,g14627);
  AN2 AND2_1747(g27697,g25785,g23649);
  AN2 AND2_1748(g18582,g2922,g16349);
  AN2 AND2_1749(g27995,g26809,g23985);
  AN2 AND2_1750(g31654,g29325,g13062);
  AN2 AND2_1751(g30576,g18898,g29800);
  AN2 AND2_1752(g22127,g6625,g19277);
  AN2 AND2_1753(g34585,g24705,g34316);
  AN2 AND2_1754(g34484,g34407,g18939);
  AN2 AND2_1755(g18310,g1333,g16931);
  AN2 AND2_1756(g29601,g1890,g28955);
  AN2 AND2_1757(g31936,g31213,g24005);
  AN2 AND2_1758(g33417,g32371,g21424);
  AN4 AND4_114(I31327,g32928,g32929,g32930,g32931);
  AN2 AND2_1759(g21789,g3451,g20391);
  AN2 AND2_1760(g26799,g25247,g21068);
  AN2 AND2_1761(g29975,g28986,g10420);
  AN2 AND2_1762(g34554,g34347,g20495);
  AN2 AND2_1763(g18627,g15093,g17093);
  AN2 AND2_1764(g15863,g13762,g13223);
  AN2 AND2_1765(g18379,g1906,g15171);
  AN2 AND2_1766(g30200,g28665,g23862);
  AN2 AND2_1767(g21788,g3401,g20391);
  AN2 AND2_1768(g33334,g32219,g20613);
  AN2 AND2_1769(g18112,g182,g17015);
  AN2 AND2_1770(g16422,g8216,g13627);
  AN2 AND2_1771(g23724,g14767,g21123);
  AN2 AND2_1772(g25852,g4593,g24411);
  AN2 AND2_1773(g18378,g1932,g15171);
  AN2 AND2_1774(g22103,g15164,g18833);
  AN3 AND3_110(g34115,g20516,g9104,g33750);
  AN2 AND2_1775(g21829,g3770,g20453);
  AN2 AND2_1776(g29937,g13044,g29196);
  AN2 AND2_1777(g14220,g8612,g11820);
  AN2 AND2_1778(g21920,g5062,g21468);
  AN2 AND2_1779(g23920,g4135,g19549);
  AN2 AND2_1780(g22095,g6428,g18833);
  AN2 AND2_1781(g16208,g3965,g14085);
  AN2 AND2_1782(g25963,g1657,g24978);
  AN2 AND2_1783(g28318,g27233,g19770);
  AN2 AND2_1784(g18386,g1964,g15171);
  AN2 AND2_1785(g30921,g29900,g24789);
  AN2 AND2_1786(g28227,g9397,g27583);
  AN2 AND2_1787(g21828,g3767,g20453);
  AN2 AND2_1788(g15703,g452,g13437);
  AN2 AND2_1789(g17784,g1152,g13215);
  AN2 AND2_1790(g23828,g9104,g19128);
  AN2 AND2_1791(g18603,g3119,g16987);
  AN2 AND2_1792(g21946,g5252,g18997);
  AN2 AND2_1793(g18742,g5120,g17847);
  AN4 AND4_115(g27445,g8038,g26314,g9187,g504);
  AN2 AND2_1794(g33423,g32225,g29657);
  AN2 AND2_1795(g29884,g2555,g29153);
  AN2 AND2_1796(g23121,g19128,g9104);
  AN2 AND2_1797(g24229,g896,g22594);
  AN2 AND2_1798(g34745,g34669,g19482);
  AN2 AND2_1799(g27316,g2407,g26710);
  AN2 AND2_1800(g24228,g862,g22594);
  AN2 AND2_1801(g18681,g4653,g15885);
  AN4 AND4_116(I31091,g29385,g32586,g32587,g32588);
  AN2 AND2_1802(g24011,g7939,g19524);
  AN2 AND2_1803(g32326,g31317,g23539);
  AN2 AND2_1804(g29666,g28980,g22498);
  AN2 AND2_1805(g17181,g1945,g13014);
  AN2 AND2_1806(g16614,g5945,g14933);
  AN2 AND2_1807(g17671,g7685,g13485);
  AN2 AND2_1808(g29363,g8458,g28444);
  AN2 AND2_1809(g23682,g16970,g20874);
  AN2 AND2_1810(g18802,g6195,g15348);
  AN2 AND2_1811(g18429,g2193,g18008);
  AN2 AND2_1812(g32040,g14122,g31243);
  AN2 AND2_1813(g24716,g15935,g23004);
  AN4 AND4_117(I24680,g24029,g24030,g24031,g24032);
  AN2 AND2_1814(g33909,g33131,g10708);
  AN2 AND2_1815(g34184,g33698,g24388);
  AN2 AND2_1816(g18730,g4950,g16861);
  AN2 AND2_1817(g15821,g3598,g14110);
  AN2 AND2_1818(g27988,g26781,g23941);
  AN2 AND2_1819(g18793,g6159,g15348);
  AN2 AND2_1820(g18428,g2169,g18008);
  AN2 AND2_1821(g24582,g5808,g23402);
  AN2 AND2_1822(g33908,g33092,g18935);
  AN3 AND3_111(g28281,g7362,g1936,g27440);
  AN2 AND2_1823(g16593,g5599,g14885);
  AN2 AND2_1824(g12924,g1570,g10980);
  AN2 AND2_1825(g27432,g26519,g17582);
  AN2 AND2_1826(g13020,g401,g11048);
  AN2 AND2_1827(g18765,g5489,g17929);
  AN2 AND2_1828(g28301,g27224,g19750);
  AN2 AND2_1829(g24310,g4495,g22228);
  AN2 AND2_1830(g16122,g9491,g14291);
  AN2 AND2_1831(g18690,g15130,g16053);
  AN4 AND4_118(g28739,g21434,g26424,g25274,g27395);
  AN2 AND2_1832(g18549,g2799,g15277);
  AN2 AND2_1833(g11046,g9889,g6120);
  AN2 AND2_1834(g25921,g24936,g9664);
  AN2 AND2_1835(g13046,g6870,g11270);
  AN2 AND2_1836(g26207,g2638,g25170);
  AN2 AND2_1837(g24627,g22763,g19679);
  AN2 AND2_1838(g29580,g28519,g14186);
  AN2 AND2_1839(g21760,g3207,g20785);
  AN2 AND2_1840(g20112,g13540,g16661);
  AN2 AND2_1841(g31242,g29373,g25409);
  AN2 AND2_1842(g22089,g6311,g19210);
  AN2 AND2_1843(g27461,g26576,g17611);
  AN2 AND2_1844(g33242,g32123,g19931);
  AN2 AND2_1845(g18548,g2807,g15277);
  AN2 AND2_1846(g15873,g3550,g14072);
  AN2 AND2_1847(g28645,g27556,g20599);
  AN4 AND4_119(I31192,g32733,g32734,g32735,g32736);
  AN2 AND2_1848(g27342,g12592,g26792);
  AN2 AND2_1849(g24378,g3106,g22718);
  AN2 AND2_1850(g16641,g6613,g14782);
  AN2 AND2_1851(g27145,g14121,g26382);
  AN2 AND2_1852(g22088,g6307,g19210);
  AN2 AND2_1853(g18504,g2579,g15509);
  AN2 AND2_1854(g22024,g5897,g19147);
  AN2 AND2_1855(g31123,g1834,g29994);
  AN2 AND2_1856(g32183,g2795,g31653);
  AN2 AND2_1857(g19266,g246,g16214);
  AN2 AND2_1858(g33814,g33098,g28144);
  AN2 AND2_1859(g28290,g23780,g27759);
  AN2 AND2_1860(g32397,g31068,g15830);
  AN2 AND2_1861(g13282,g3546,g11480);
  AN2 AND2_1862(g27650,g26519,g15479);
  AN4 AND4_120(g29110,g27187,g12687,g20751,I27429);
  AN2 AND2_1863(g25973,g2342,g24994);
  AN2 AND2_1864(g18317,g12846,g17873);
  AN2 AND2_1865(g33807,g33112,g25452);
  AN2 AND2_1866(g31974,g31760,g22176);
  AN2 AND2_1867(g29321,g29033,g22148);
  AN2 AND2_1868(g33639,g33386,g18829);
  AN4 AND4_121(g26241,g24688,g10678,g8778,g10627);
  AN2 AND2_1869(g34214,g33772,g22689);
  AN2 AND2_1870(g29531,g1664,g28559);
  AN2 AND2_1871(g31230,g30285,g20751);
  AN2 AND2_1872(g18129,g518,g16971);
  AN2 AND2_1873(g30207,g28680,g23874);
  AN2 AND2_1874(g16635,g5607,g14959);
  AN2 AND2_1875(g27696,g25800,g23647);
  AN2 AND2_1876(g34329,g14511,g34181);
  AN2 AND2_1877(g27330,g2541,g26744);
  AN2 AND2_1878(g27393,g26099,g20066);
  AN2 AND2_1879(g28427,g27258,g20008);
  AN2 AND2_1880(g24681,g16653,g22988);
  AN2 AND2_1881(g29178,g27163,g12687);
  AN2 AND2_1882(g29740,g2648,g29154);
  AN2 AND2_1883(g30005,g28230,g24394);
  AN2 AND2_1884(g22126,g6621,g19277);
  AN2 AND2_1885(g18128,g504,g16971);
  AN2 AND2_1886(g21927,g5164,g18997);
  AN2 AND2_1887(g26100,g1677,g25097);
  AN2 AND2_1888(g19588,g3849,g16853);
  AN2 AND2_1889(g33416,g32370,g21423);
  AN2 AND2_1890(g29685,g2084,g28711);
  AN4 AND4_122(I31326,g30735,g31853,g32926,g32927);
  AN2 AND2_1891(g18245,g1193,g16431);
  AN2 AND2_1892(g27132,g26055,g16589);
  AN2 AND2_1893(g34538,g34330,g20054);
  AN2 AND2_1894(g18626,g3498,g17062);
  AN2 AND2_1895(g15913,g3933,g14021);
  AN2 AND2_1896(g24730,g6177,g23699);
  AN2 AND2_1897(g31992,g31773,g22213);
  AN2 AND2_1898(g18323,g1632,g17873);
  AN2 AND2_1899(g33841,g33254,g20268);
  AN2 AND2_1900(g18299,g1526,g16489);
  AN2 AND2_1901(g18533,g2729,g15277);
  AN2 AND2_1902(g28547,g6821,g27091);
  AN3 AND3_112(g33510,g32816,I31246,I31247);
  AN2 AND2_1903(g24765,g17699,g22498);
  AN2 AND2_1904(g18298,g15073,g16489);
  AN3 AND3_113(g27161,g26166,g8241,g1783);
  AN2 AND2_1905(g30241,g28729,g23926);
  AN4 AND4_123(I31252,g32819,g32820,g32821,g32822);
  AN2 AND2_1906(g31579,g19128,g29814);
  AN2 AND2_1907(g18775,g7028,g15615);
  AN2 AND2_1908(g24549,g23162,g20887);
  AN2 AND2_1909(g28226,g27825,g26667);
  AN2 AND2_1910(g21755,g3203,g20785);
  AN2 AND2_1911(g29334,g29148,g18908);
  AN2 AND2_1912(g16474,g8280,g13666);
  AN2 AND2_1913(g23755,g14821,g21204);
  AN2 AND2_1914(g27259,g26755,g26725);
  AN2 AND2_1915(g19749,g732,g16646);
  AN2 AND2_1916(g32047,g27248,g31070);
  AN2 AND2_1917(g33835,g4340,g33413);
  AN2 AND2_1918(g9968,g1339,g1500);
  AN2 AND2_1919(g21770,g3251,g20785);
  AN2 AND2_1920(g32205,g30922,g28463);
  AN2 AND2_1921(g21981,g5543,g19074);
  AN2 AND2_1922(g22060,g6151,g21611);
  AN2 AND2_1923(g10902,g7858,g1129);
  AN2 AND2_1924(g18737,g4975,g16826);
  AN2 AND2_1925(g27087,g13872,g26284);
  AN2 AND2_1926(g28572,g27829,g15669);
  AN2 AND2_1927(g12259,g9480,g640);
  AN2 AND2_1928(g24504,g22226,g19410);
  AN2 AND2_1929(g32311,g31295,g20582);
  AN2 AND2_1930(g25207,g22513,g10621);
  AN2 AND2_1931(g29762,g28298,g10233);
  AN2 AND2_1932(g18232,g1124,g16326);
  AN2 AND2_1933(g34771,g34693,g20147);
  AN2 AND2_1934(g29964,g2008,g28830);
  AN2 AND2_1935(g16537,g5937,g14855);
  AN2 AND2_1936(g11027,g5097,g9724);
  AN2 AND2_1937(g30235,g28723,g23915);
  AN3 AND3_114(I18713,g13156,g6767,g6756);
  AN3 AND3_115(g25328,g5022,g23764,I24505);
  AN2 AND2_1938(g11890,g7499,g9155);
  AN2 AND2_1939(g24317,g4534,g22228);
  AN2 AND2_1940(g15797,g3909,g14139);
  AN2 AND2_1941(g18697,g4749,g16777);
  AN2 AND2_1942(g27043,g26335,g8632);
  AN2 AND2_1943(g32051,g31506,g10831);
  AN4 AND4_124(g16283,g11547,g11592,g6789,I17606);
  AN2 AND2_1944(g29587,g2181,g28935);
  AN4 AND4_125(I31062,g32545,g32546,g32547,g32548);
  AN2 AND2_1945(g18261,g1256,g16000);
  AN2 AND2_1946(g21767,g3239,g20785);
  AN2 AND2_1947(g21794,g15094,g20924);
  AN2 AND2_1948(g21845,g3881,g21070);
  AN2 AND2_1949(g12043,g1345,g7601);
  AN2 AND2_1950(g16303,g4527,g12921);
  AN2 AND2_1951(g10290,g4358,g4349);
  AN2 AND2_1952(g24002,g19613,g10971);
  AN2 AND2_1953(g21990,g5591,g19074);
  AN2 AND2_1954(g11003,g7880,g1300);
  AN2 AND2_1955(g18512,g2619,g15509);
  AN2 AND2_1956(g23990,g19610,g10951);
  AN4 AND4_126(I27524,g28037,g24114,g24115,g24116);
  AN2 AND2_1957(g33720,g33161,g19439);
  AN3 AND3_116(g19560,g15832,g1157,g10893);
  AN2 AND2_1958(g29909,g28435,g23388);
  AN4 AND4_127(g27602,g23032,g26244,g26424,g24966);
  AN2 AND2_1959(g31275,g30147,g27800);
  AN2 AND2_1960(g34515,g34288,g19491);
  AN2 AND2_1961(g34414,g34206,g21457);
  AN4 AND4_128(g28889,g17292,g25169,g26424,g27395);
  AN2 AND2_1962(g31746,g30093,g23905);
  AN2 AND2_1963(g27375,g26519,g17479);
  AN2 AND2_1964(g26206,g2523,g25495);
  AN2 AND2_1965(g31493,g29791,g23434);
  AN2 AND2_1966(g32350,g2697,g31710);
  AN2 AND2_1967(g21719,g358,g21037);
  AN3 AND3_117(g33493,g32693,I31161,I31162);
  AN2 AND2_1968(g24323,g4546,g22228);
  AN2 AND2_1969(g24299,g4456,g22550);
  AN2 AND2_1970(g13778,g4540,g10597);
  AN2 AND2_1971(g13081,g8626,g11122);
  AN2 AND2_1972(g29569,g29028,g22498);
  AN2 AND2_1973(g21718,g370,g21037);
  AN3 AND3_118(g33465,g32491,I31021,I31022);
  AN2 AND2_1974(g31237,g29366,g25325);
  AN3 AND3_119(g10632,g7475,g7441,g890);
  AN2 AND2_1975(g24298,g4392,g22550);
  AN2 AND2_1976(g33237,g32394,g25198);
  AN2 AND2_1977(g32152,g31631,g29998);
  AN2 AND2_1978(g18445,g2273,g18008);
  AN2 AND2_1979(g24775,g17594,g22498);
  AN2 AND2_1980(g29568,g2571,g28950);
  AN2 AND2_1981(g29747,g28286,g23196);
  AN2 AND2_1982(g32396,g4698,g30983);
  AN2 AND2_1983(g33340,g32222,g20639);
  AN2 AND2_1984(g21832,g3787,g20453);
  AN2 AND2_1985(g18499,g2476,g15426);
  AN2 AND2_1986(g18316,g1564,g16931);
  AN2 AND2_1987(g33684,g33139,g13565);
  AN2 AND2_1988(g16840,g5467,g14262);
  AN2 AND2_1989(g31142,g2527,g30039);
  AN2 AND2_1990(g22055,g6128,g21611);
  AN2 AND2_1991(g18498,g2547,g15426);
  AN2 AND2_1992(g32413,g31121,g19518);
  AN2 AND2_1993(g19693,g6181,g17087);
  AN2 AND2_1994(g22111,g6549,g19277);
  AN4 AND4_129(I31047,g32524,g32525,g32526,g32527);
  AN2 AND2_1995(g21861,g3949,g21070);
  AN2 AND2_1996(g34584,g24653,g34315);
  AN2 AND2_1997(g22070,g6243,g19210);
  AN2 AND2_1998(g13998,g6589,g12629);
  AN2 AND2_1999(g31517,g29849,g23482);
  AN2 AND2_2000(g26345,g13051,g25505);
  AN2 AND2_2001(g28426,g27257,g20006);
  AN3 AND3_120(g33517,g32867,I31281,I31282);
  AN2 AND2_2002(g29751,g28297,g23216);
  AN2 AND2_2003(g29807,g28359,g23272);
  AN4 AND4_130(I31311,g30673,g31851,g32903,g32904);
  AN2 AND2_2004(g29772,g28323,g23243);
  AN2 AND2_2005(g22590,g19274,g19452);
  AN2 AND2_2006(g16192,g6191,g14321);
  AN2 AND2_2007(g26849,g2994,g24527);
  AN2 AND2_2008(g29974,g29173,g12914);
  AN2 AND2_2009(g15711,g460,g13437);
  AN2 AND2_2010(g18611,g15090,g17200);
  AN2 AND2_2011(g27459,g26549,g17609);
  AN2 AND2_2012(g21926,g15147,g18997);
  AN2 AND2_2013(g18722,g4917,g16077);
  AN2 AND2_2014(g26399,g15572,g25566);
  AN3 AND3_121(g25414,g5406,g22194,I24549);
  AN2 AND2_2015(g25991,g2060,g25023);
  AN2 AND2_2016(g23389,g9072,g19757);
  AN2 AND2_2017(g29639,g28510,g11618);
  AN2 AND2_2018(g15109,g4269,g14454);
  AN2 AND2_2019(g26848,g2950,g24526);
  AN3 AND3_122(I16646,g10160,g12413,g12343);
  AN2 AND2_2020(g26398,g24946,g10474);
  AN3 AND3_123(g22384,g9354,g9285,g20784);
  AN2 AND2_2021(g18432,g2223,g18008);
  AN4 AND4_131(I24705,g24064,g24065,g24066,g24067);
  AN2 AND2_2022(g29638,g2583,g29025);
  AN4 AND4_132(I31051,g31376,g31804,g32529,g32530);
  AN2 AND2_2023(g21701,g153,g20283);
  AN4 AND4_133(I31072,g32559,g32560,g32561,g32562);
  AN2 AND2_2024(g18271,g1296,g16031);
  AN2 AND2_2025(g30082,g29181,g12752);
  AN2 AND2_2026(g34114,g33920,g23742);
  AN2 AND2_2027(g15108,g4264,g14454);
  AN2 AND2_2028(g21777,g3380,g20391);
  AN2 AND2_2029(g34758,g34683,g19657);
  AN2 AND2_2030(g26652,g10799,g24426);
  AN2 AND2_2031(g31130,g12191,g30019);
  AN2 AND2_2032(g22067,g6215,g19210);
  AN2 AND2_2033(g22094,g6398,g18833);
  AN2 AND2_2034(g34082,g33709,g19554);
  AN2 AND2_2035(g30107,g28560,g20909);
  AN2 AND2_2036(g21251,g13969,g17470);
  AN4 AND4_134(I24679,g19968,g24026,g24027,g24028);
  AN2 AND2_2037(g33362,g32259,g20914);
  AN2 AND2_2038(g11449,g6052,g7175);
  AN2 AND2_2039(g27545,g26519,g17756);
  AN2 AND2_2040(g16483,g5224,g14915);
  AN2 AND2_2041(g18753,g15148,g15595);
  AN2 AND2_2042(g18461,g2307,g15224);
  AN2 AND2_2043(g31523,g7528,g29333);
  AN2 AND2_2044(g32020,g4157,g30937);
  AN2 AND2_2045(g18342,g1592,g17873);
  AN3 AND3_124(g33523,g32909,I31311,I31312);
  AN2 AND2_2046(g29841,g28371,g23283);
  AN2 AND2_2047(g19914,g2815,g15853);
  AN2 AND2_2048(g29992,g29012,g10490);
  AN2 AND2_2049(g27599,g26337,g20033);
  AN2 AND2_2050(g34744,g34668,g19481);
  AN2 AND2_2051(g18145,g582,g17533);
  AN2 AND2_2052(g29510,g28856,g22342);
  AN2 AND2_2053(g32046,g10925,g30735);
  AN2 AND2_2054(g18199,g832,g17821);
  AN2 AND2_2055(g22019,g5857,g19147);
  AN2 AND2_2056(g27598,g25899,g10475);
  AN2 AND2_2057(g18650,g6928,g17271);
  AN2 AND2_2058(g18736,g4991,g16826);
  AN2 AND2_2059(g27086,g25836,g22495);
  AN2 AND2_2060(g31475,g29756,g23406);
  AN2 AND2_2061(g29579,g28457,g7964);
  AN2 AND2_2062(g17150,g8579,g12995);
  AN3 AND3_125(I24030,g8390,g8016,g3396);
  AN3 AND3_126(g33475,g32563,I31071,I31072);
  AN2 AND2_2063(g16536,g5917,g14996);
  AN2 AND2_2064(g18198,g15059,g17821);
  AN2 AND2_2065(g22018,g15157,g19147);
  AN2 AND2_2066(g18529,g2712,g15277);
  AN2 AND2_2067(g21997,g5619,g19074);
  AN2 AND2_2068(g32113,g31601,g29925);
  AN2 AND2_2069(g34398,g7684,g34070);
  AN4 AND4_135(I31152,g32675,g32676,g32677,g32678);
  AN2 AND2_2070(g33727,g33115,g19499);
  AN2 AND2_2071(g24499,g22217,g19394);
  AN2 AND2_2072(g29578,g2491,g28606);
  AN2 AND2_2073(g33863,g33273,g20505);
  AN2 AND2_2074(g19594,g11913,g17268);
  AN2 AND2_2075(g29835,g28326,g24866);
  AN2 AND2_2076(g34141,g33932,g23828);
  AN2 AND2_2077(g16702,g5615,g14691);
  AN2 AND2_2078(g24316,g4527,g22228);
  AN2 AND2_2079(g31222,g2643,g30113);
  AN2 AND2_2080(g32282,g31258,g20503);
  AN4 AND4_136(g27817,g22498,g25245,g26424,g26236);
  AN2 AND2_2081(g15796,g3586,g14015);
  AN2 AND2_2082(g18696,g4741,g16053);
  AN2 AND2_2083(g18330,g1668,g17873);
  AN2 AND2_2084(g32302,g31279,g23485);
  AN2 AND2_2085(g18393,g1917,g15171);
  AN2 AND2_2086(g24498,g14036,g23850);
  AN2 AND2_2087(g29586,g1886,g28927);
  AN2 AND2_2088(g16621,g8278,g13821);
  AN2 AND2_2089(g12817,g1351,g7601);
  AN2 AND2_2090(g21766,g3235,g20785);
  AN2 AND2_2091(g26833,g2852,g24509);
  AN2 AND2_2092(g26049,g9621,g25046);
  AN2 AND2_2093(g30263,g28773,g23962);
  AN2 AND2_2094(g32105,g4922,g30673);
  AN2 AND2_2095(g28658,g27563,g20611);
  AN2 AND2_2096(g18764,g5485,g17929);
  AN4 AND4_137(g20056,g16291,g9007,g8954,g8903);
  AN2 AND2_2097(g18365,g1848,g17955);
  AN2 AND2_2098(g27158,g26609,g16645);
  AN2 AND2_2099(g21871,g4108,g19801);
  AN2 AND2_2100(g25107,g17643,g23508);
  AN3 AND3_127(g22457,g7753,g7717,g21288);
  AN2 AND2_2101(g15840,g3949,g14142);
  AN2 AND2_2102(g18132,g513,g16971);
  AN2 AND2_2103(g26048,g5853,g25044);
  AN2 AND2_2104(g28339,g9946,g27693);
  AN2 AND2_2105(g30135,g28592,g21180);
  AN2 AND2_2106(g24722,g17618,g22417);
  AN2 AND2_2107(g34135,g33926,g23802);
  AN3 AND3_128(I18782,g13156,g11450,g6756);
  AN2 AND2_2108(g7948,g1548,g1430);
  AN2 AND2_2109(g29615,g1844,g29049);
  AN2 AND2_2110(g16673,g6617,g14822);
  AN2 AND2_2111(g18161,g691,g17433);
  AN2 AND2_2112(g34962,g34945,g23020);
  AN2 AND2_2113(g19637,g5142,g16958);
  AN2 AND2_2114(g26613,g1361,g24518);
  AN2 AND2_2115(g18709,g59,g17302);
  AN2 AND2_2116(g22001,g5731,g21562);
  AN2 AND2_2117(g22077,g6263,g19210);
  AN2 AND2_2118(g25848,g25539,g18977);
  AN2 AND2_2119(g14190,g859,g10632);
  AN2 AND2_2120(g27336,g2675,g26777);
  AN2 AND2_2121(g30049,g13114,g28167);
  AN2 AND2_2122(g18259,g15068,g16000);
  AN2 AND2_2123(g29746,g28279,g20037);
  AN2 AND2_2124(g34500,g34276,g30568);
  AN2 AND2_2125(g18225,g1041,g16100);
  AN2 AND2_2126(g33351,g32236,g20707);
  AN2 AND2_2127(g33372,g32285,g21183);
  AN2 AND2_2128(g18708,g4818,g16782);
  AN2 AND2_2129(g28197,g27647,g11344);
  AN2 AND2_2130(g25804,g8069,g24587);
  AN2 AND2_2131(g18471,g2407,g15224);
  AN2 AND2_2132(g33821,g33238,g20153);
  AN2 AND2_2133(g26273,g2122,g25389);
  AN2 AND2_2134(g30048,g29193,g12945);
  AN2 AND2_2135(g22689,g18918,g9104);
  AN2 AND2_2136(g18258,g1221,g16897);
  AN2 AND2_2137(g16634,g5264,g14953);
  AN2 AND2_2138(g20887,g16282,g4864);
  AN2 AND2_2139(g23451,g13805,g20510);
  AN2 AND2_2140(g24199,g355,g22722);
  AN2 AND2_2141(g24650,g22641,g19718);
  AN2 AND2_2142(g23220,g19417,g20067);
  AN3 AND3_129(g24887,g3712,g23239,I24054);
  AN2 AND2_2143(g30004,g28521,g25837);
  AN4 AND4_138(I31046,g29385,g32521,g32522,g32523);
  AN2 AND2_2144(g22624,g19344,g19471);
  AN2 AND2_2145(g21911,g5046,g21468);
  AN2 AND2_2146(g30221,g28700,g23893);
  AN2 AND2_2147(g31790,g21299,g29385);
  AN2 AND2_2148(g33264,g31965,g21306);
  AN2 AND2_2149(g31516,g29848,g23476);
  AN2 AND2_2150(g24198,g351,g22722);
  AN2 AND2_2151(g33790,g33108,g20643);
  AN3 AND3_130(g33516,g32860,I31276,I31277);
  AN2 AND2_2152(g29806,g28358,g23271);
  AN2 AND2_2153(g29684,g1982,g29085);
  AN2 AND2_2154(g18244,g1171,g16431);
  AN2 AND2_2155(g26234,g2657,g25514);
  AN2 AND2_2156(g22102,g6479,g18833);
  AN3 AND3_131(g24843,g3010,g23211,I24015);
  AN2 AND2_2157(g33873,g33291,g20549);
  AN2 AND2_2158(g24330,g18661,g22228);
  AN2 AND2_2159(g22157,g14608,g18892);
  AN2 AND2_2160(g24393,g3808,g22844);
  AN3 AND3_132(I24075,g3736,g3742,g8553);
  AN4 AND4_139(I31282,g32863,g32864,g32865,g32866);
  AN2 AND2_2161(g25962,g9258,g24971);
  AN4 AND4_140(g16213,g6772,g6782,g11640,I17552);
  AN2 AND2_2162(g24764,g17570,g22472);
  AN2 AND2_2163(g29517,g1870,g28827);
  AN4 AND4_141(I31302,g32891,g32892,g32893,g32894);
  AN4 AND4_142(I31357,g32970,g32971,g32972,g32973);
  AN2 AND2_2164(g21776,g3376,g20391);
  AN2 AND2_2165(g21785,g3431,g20391);
  AN4 AND4_143(I27519,g28036,g24107,g24108,g24109);
  AN2 AND2_2166(g18602,g3115,g16987);
  AN2 AND2_2167(g18810,g6505,g15483);
  AN2 AND2_2168(g15757,g3207,g14066);
  AN2 AND2_2169(g18657,g4308,g17128);
  AN2 AND2_2170(g22066,g6209,g19210);
  AN2 AND2_2171(g18774,g5698,g15615);
  AN2 AND2_2172(g7918,g1205,g1087);
  AN2 AND2_2173(g18375,g1902,g15171);
  AN2 AND2_2174(g31209,g2084,g30097);
  AN2 AND2_2175(g33422,g32375,g21456);
  AN2 AND2_2176(g34106,g33917,g23675);
  AN2 AND2_2177(g32248,g31616,g30299);
  AN2 AND2_2178(g21754,g3195,g20785);
  AN4 AND4_144(I27518,g20720,g24104,g24105,g24106);
  AN2 AND2_2179(g10625,g3431,g7926);
  AN2 AND2_2180(g27309,g26603,g23057);
  AN2 AND2_2181(g23754,g14816,g21189);
  AN2 AND2_2182(g28714,g27591,g20711);
  AN3 AND3_133(g16047,g13322,g1500,g10699);
  AN2 AND2_2183(g25833,g8228,g24626);
  AN2 AND2_2184(g14126,g881,g10632);
  AN4 AND4_145(g16205,g11547,g6782,g11640,I17542);
  AN2 AND2_2185(g27288,g26515,g23013);
  AN2 AND2_2186(g28315,g27232,g19769);
  AN2 AND2_2187(g33834,g33095,g29172);
  AN2 AND2_2188(g31208,g30262,g25188);
  AN2 AND2_2189(g32204,g4245,g31327);
  AN2 AND2_2190(g21859,g3941,g21070);
  AN2 AND2_2191(g21825,g3736,g20453);
  AN2 AND2_2192(g21950,g5268,g18997);
  AN2 AND2_2193(g26514,g7400,g25564);
  AN2 AND2_2194(g22876,g20136,g9104);
  AN2 AND2_2195(g18337,g1706,g17873);
  AN2 AND2_2196(g28202,g27659,g11413);
  AN2 AND2_2197(g30033,g29189,g12937);
  AN2 AND2_2198(g28257,g27179,g19686);
  AN2 AND2_2199(g21858,g3937,g21070);
  AN2 AND2_2200(g29362,g27379,g28307);
  AN2 AND2_2201(g18171,g728,g17433);
  AN2 AND2_2202(g30234,g28721,g23914);
  AN2 AND2_2203(g34371,g7450,g34044);
  AN2 AND2_2204(g24709,g16690,g23000);
  AN2 AND2_2205(g31542,g19050,g29814);
  AN2 AND2_2206(g31021,g26025,g29814);
  AN2 AND2_2207(g29523,g28930,g22417);
  AN2 AND2_2208(g23151,g18994,g7162);
  AN2 AND2_2209(g28111,g27343,g22716);
  AN2 AND2_2210(g14296,g2638,g11897);
  AN2 AND2_2211(g21996,g5615,g19074);
  AN2 AND2_2212(g24225,g246,g22594);
  AN2 AND2_2213(g15673,g182,g13437);
  AN2 AND2_2214(g18792,g7051,g15634);
  AN2 AND2_2215(g15847,g3191,g14005);
  AN2 AND2_2216(g23996,g19596,g10951);
  AN2 AND2_2217(g24708,g16474,g22998);
  AN2 AND2_2218(g14644,g10610,g10605);
  AN3 AND3_134(g33913,g23088,g33204,g9104);
  AN2 AND2_2219(g16592,g5579,g14688);
  AN2 AND2_2220(g21844,g3873,g21070);
  AN2 AND2_2221(g21394,g13335,g15799);
  AN2 AND2_2222(g32356,g2704,g31710);
  AN2 AND2_2223(g29475,g14033,g28500);
  AN2 AND2_2224(g18459,g2331,g15224);
  AN2 AND2_2225(g18425,g2161,g18008);
  AN2 AND2_2226(g33905,g33089,g15574);
  AN2 AND2_2227(g33073,g32386,g18828);
  AN2 AND2_2228(g12687,g9024,g8977);
  AN2 AND2_2229(g25106,g17391,g23506);
  AN2 AND2_2230(g26541,g319,g24375);
  AN2 AND2_2231(g34514,g34286,g19480);
  AN2 AND2_2232(g15851,g3953,g14157);
  AN2 AND2_2233(g15872,g9095,g14234);
  AN2 AND2_2234(g18458,g2357,g15224);
  AN2 AND2_2235(g19139,g452,g16195);
  AN2 AND2_2236(g27374,g26519,g17478);
  AN3 AND3_135(g33530,g32960,I31346,I31347);
  AN2 AND2_2237(g21420,g16093,g13596);
  AN2 AND2_2238(g34507,g34280,g19454);
  AN2 AND2_2239(g31122,g12144,g29993);
  AN2 AND2_2240(g32182,g31753,g27937);
  AN4 AND4_146(g20069,g16312,g9051,g9011,g8955);
  AN2 AND2_2241(g33122,g8859,g32192);
  AN2 AND2_2242(g8530,g2902,g2907);
  AN4 AND4_147(I31027,g32494,g32495,g32496,g32497);
  AN3 AND3_136(I24524,g5041,g5046,g9716);
  AN3 AND3_137(g33464,g32484,I31016,I31017);
  AN3 AND3_138(I16129,g8728,g11443,g11411);
  AN2 AND2_2243(g20602,g10803,g15580);
  AN4 AND4_148(g28150,g10862,g11834,g11283,g27187);
  AN3 AND3_139(g16846,g14034,g12591,g11185);
  AN2 AND2_2244(g18545,g2783,g15277);
  AN2 AND2_2245(g25951,g24500,g19565);
  AN2 AND2_2246(g26325,g12644,g25370);
  AN2 AND2_2247(g24602,g16507,g22854);
  AN2 AND2_2248(g25972,g2217,g24993);
  AN2 AND2_2249(g18444,g2269,g18008);
  AN2 AND2_2250(g25033,g17500,g23433);
  AN3 AND3_140(g25371,g5062,g22173,I24524);
  AN2 AND2_2251(g20375,g671,g16846);
  AN2 AND2_2252(g24657,g22644,g19730);
  AN2 AND2_2253(g24774,g718,g23614);
  AN2 AND2_2254(g16731,g7153,g12941);
  AN2 AND2_2255(g26829,g2844,g24505);
  AN2 AND2_2256(g27669,g26840,g13278);
  AN2 AND2_2257(g17480,g9683,g14433);
  AN2 AND2_2258(g19333,g464,g16223);
  AN2 AND2_2259(g29347,g29176,g22201);
  AN2 AND2_2260(g18599,g2955,g16349);
  AN2 AND2_2261(g22307,g20027,g21163);
  AN2 AND2_2262(g22076,g6255,g19210);
  AN2 AND2_2263(g22085,g6295,g19210);
  AN2 AND2_2264(g26358,g19522,g25528);
  AN3 AND3_141(I27349,g25534,g26424,g22698);
  AN2 AND2_2265(g23025,g16021,g19798);
  AN2 AND2_2266(g27260,g26766,g26737);
  AN2 AND2_2267(g32331,g31322,g20637);
  AN2 AND2_2268(g31292,g29735,g23338);
  AN2 AND2_2269(g26828,g24919,g15756);
  AN2 AND2_2270(g27668,g1367,g25917);
  AN2 AND2_2271(g23540,g16866,g20622);
  AN2 AND2_2272(g18598,g3003,g16349);
  AN2 AND2_2273(g22054,g6120,g21611);
  AN2 AND2_2274(g28695,g27580,g20666);
  AN2 AND2_2275(g31153,g12336,g30068);
  AN2 AND2_2276(g27392,g26576,g17507);
  AN2 AND2_2277(g29600,g1840,g29049);
  AN2 AND2_2278(g26121,g6167,g25111);
  AN2 AND2_2279(g20171,g16479,g10476);
  AN2 AND2_2280(g34541,g34331,g20087);
  AN2 AND2_2281(g17307,g9498,g14343);
  AN2 AND2_2282(g15574,g4311,g13202);
  AN2 AND2_2283(g33409,g32359,g21408);
  AN3 AND3_142(I24616,g6082,g6088,g9946);
  AN2 AND2_2284(g29952,g23576,g28939);
  AN2 AND2_2285(g27559,g26576,g17777);
  AN2 AND2_2286(g29351,g4771,g28406);
  AN2 AND2_2287(g27525,g26576,g17720);
  AN2 AND2_2288(g27488,g26549,g17648);
  AN2 AND2_2289(g18817,g6533,g15483);
  AN2 AND2_2290(g15912,g3562,g14018);
  AN4 AND4_149(g14581,g12587,g12428,g12357,I16695);
  AN2 AND2_2291(g18322,g1608,g17873);
  AN2 AND2_2292(g33408,g32358,g21407);
  AN4 AND4_150(I31081,g30673,g31810,g32571,g32572);
  AN2 AND2_2293(g24967,g23197,g20213);
  AN2 AND2_2294(g10707,g3787,g8561);
  AN2 AND2_2295(g18159,g671,g17433);
  AN2 AND2_2296(g27558,g26576,g17776);
  AN3 AND3_143(g25507,g6098,g23844,I24616);
  AN2 AND2_2297(g22942,g9104,g20219);
  AN2 AND2_2298(g18125,g15053,g16886);
  AN2 AND2_2299(g18532,g2724,g15277);
  AN2 AND2_2300(g26291,g2681,g25439);
  AN2 AND2_2301(g30920,g29889,g21024);
  AN4 AND4_151(I24704,g21193,g24061,g24062,g24063);
  AN2 AND2_2302(g19585,g17180,g14004);
  AN2 AND2_2303(g14202,g869,g10632);
  AN2 AND2_2304(g16929,g6505,g14348);
  AN2 AND2_2305(g18158,g667,g17433);
  AN2 AND2_2306(g14257,g8612,g11878);
  AN2 AND2_2307(g21957,g5390,g21514);
  AN2 AND2_2308(g18783,g5841,g18065);
  AN2 AND2_2309(g23957,g4138,g19589);
  AN2 AND2_2310(g29516,g28895,g22369);
  AN4 AND4_152(g14496,g12411,g12244,g12197,I16618);
  AN2 AND2_2311(g22670,g20114,g9104);
  AN2 AND2_2312(g21739,g3080,g20330);
  AN4 AND4_153(I31356,g31327,g31859,g32968,g32969);
  AN2 AND2_2313(g25163,g20217,g23566);
  AN2 AND2_2314(g18561,g2841,g15277);
  AN2 AND2_2315(g18656,g15120,g17128);
  AN2 AND2_2316(g30121,g28577,g21052);
  AN2 AND2_2317(g25012,g20644,g23419);
  AN2 AND2_2318(g18353,g1772,g17955);
  AN2 AND2_2319(g18295,g1489,g16449);
  AN2 AND2_2320(g21738,g3072,g20330);
  AN3 AND3_144(g10590,g7246,g7392,I13937);
  AN2 AND2_2321(g17156,g305,g13385);
  AN2 AND2_2322(g17655,g7897,g13342);
  AN2 AND2_2323(g18680,g15128,g15885);
  AN2 AND2_2324(g18144,g590,g17533);
  AN2 AND2_2325(g18823,g6727,g15680);
  AN2 AND2_2326(g34344,g34107,g20038);
  AN2 AND2_2327(g21699,g142,g20283);
  AN2 AND2_2328(g28706,g27584,g20681);
  AN2 AND2_2329(g28597,g27515,g20508);
  AN4 AND4_154(I31182,g32719,g32720,g32721,g32722);
  AN2 AND2_2330(g18336,g1700,g17873);
  AN2 AND2_2331(g24545,g3333,g23285);
  AN3 AND3_145(g33474,g32556,I31066,I31067);
  AN2 AND2_2332(g28256,g11398,g27984);
  AN2 AND2_2333(g15820,g3578,g13955);
  AN2 AND2_2334(g28689,g27575,g20651);
  AN2 AND2_2335(g32149,g31658,g29983);
  AN2 AND2_2336(g27042,g25774,g19343);
  AN3 AND3_146(g33711,g33176,g10727,g22332);
  AN2 AND2_2337(g30173,g28118,g13082);
  AN2 AND2_2338(g34291,g34055,g19366);
  AN2 AND2_2339(g31327,g19200,g29814);
  AN2 AND2_2340(g27255,g25936,g19689);
  AN2 AND2_2341(g28280,g23761,g27724);
  AN2 AND2_2342(g22131,g6641,g19277);
  AN2 AND2_2343(g29834,g28368,g23278);
  AN2 AND2_2344(g33327,g32208,g20561);
  AN2 AND2_2345(g34173,g33679,g24368);
  AN3 AND3_147(I24064,g3385,g3391,g8492);
  AN3 AND3_148(g29208,g24138,I27538,I27539);
  AN2 AND2_2346(g25788,g8010,g24579);
  AN2 AND2_2347(g32148,g31631,g29981);
  AN2 AND2_2348(g28624,g22357,g27009);
  AN2 AND2_2349(g28300,g27771,g26605);
  AN2 AND2_2350(g27270,g26805,g26793);
  AN2 AND2_2351(g32097,g25960,g31021);
  AN4 AND4_155(I31331,g30825,g31854,g32933,g32934);
  AN2 AND2_2352(g27678,g947,g25830);
  AN2 AND2_2353(g18631,g3694,g17226);
  AN2 AND2_2354(g32104,g31616,g29906);
  AN3 AND3_149(g7520,g2704,g2697,g2689);
  AN2 AND2_2355(g18364,g1844,g17955);
  AN2 AND2_2356(g32343,g31473,g20710);
  AN2 AND2_2357(g31283,g30156,g27837);
  AN2 AND2_2358(g27460,g26549,g17610);
  AN2 AND2_2359(g27686,g1291,g25849);
  AN2 AND2_2360(g25946,g24496,g19537);
  AN2 AND2_2361(g31492,g29790,g23431);
  AN2 AND2_2362(g24817,g22929,g7235);
  AN2 AND2_2363(g30029,g29164,g12936);
  AN3 AND3_150(g33492,g32686,I31156,I31157);
  AN2 AND2_2364(g19674,g2819,g15867);
  AN2 AND2_2365(g24322,g4423,g22228);
  AN2 AND2_2366(g12939,g405,g11048);
  AN2 AND2_2367(g27030,g26343,g7947);
  AN2 AND2_2368(g20977,g10123,g17301);
  AN2 AND2_2369(g13299,g437,g11048);
  AN2 AND2_2370(g24532,g22331,g19478);
  AN2 AND2_2371(g32369,g2130,g31672);
  AN2 AND2_2372(g27267,g26026,g17124);
  AN2 AND2_2373(g27294,g9975,g26656);
  AN2 AND2_2374(g29614,g28860,g22369);
  AN2 AND2_2375(g30028,g29069,g9311);
  AN3 AND3_151(g28231,g27187,g22763,g27074);
  AN2 AND2_2376(g24977,g23209,g20232);
  AN2 AND2_2377(g34506,g8833,g34354);
  AN2 AND2_2378(g16803,g5933,g14810);
  AN2 AND2_2379(g31750,g30103,g23925);
  AN2 AND2_2380(g29607,g28509,g14208);
  AN2 AND2_2381(g18289,g1448,g16449);
  AN4 AND4_156(I31026,g31194,g31800,g32492,g32493);
  AN2 AND2_2382(g29320,g29068,g22147);
  AN2 AND2_2383(g33381,g11842,g32318);
  AN4 AND4_157(I31212,g32761,g32762,g32763,g32764);
  AN4 AND4_158(g29073,g27163,g10290,g21012,I27409);
  AN2 AND2_2384(g12065,g9557,g9805);
  AN2 AND2_2385(g18309,g1339,g16931);
  AN2 AND2_2386(g29530,g1612,g28820);
  AN2 AND2_2387(g24656,g11736,g22926);
  AN2 AND2_2388(g29593,g28470,g7985);
  AN2 AND2_2389(g33091,g32392,g18897);
  AN2 AND2_2390(g18288,g1454,g16449);
  AN2 AND2_2391(g18224,g1036,g16100);
  AN2 AND2_2392(g21715,g160,g20283);
  AN2 AND2_2393(g22039,g5949,g19147);
  AN2 AND2_2394(g29346,g4894,g28381);
  AN2 AND2_2395(g25173,g12234,g23589);
  AN2 AND2_2396(g24295,g4434,g22550);
  AN2 AND2_2397(g18571,g2856,g16349);
  AN2 AND2_2398(g18308,g6832,g16931);
  AN2 AND2_2399(g24680,g16422,g22986);
  AN2 AND2_2400(g27219,g26026,g16742);
  AN2 AND2_2401(g32412,g4765,g30998);
  AN2 AND2_2402(g24144,g17727,g21660);
  AN2 AND2_2403(g33796,g33117,g25267);
  AN2 AND2_2404(g19692,g12066,g17086);
  AN3 AND3_152(I24555,g9559,g9809,g6093);
  AN2 AND2_2405(g29565,g1932,g28590);
  AN2 AND2_2406(g26604,g13248,g25051);
  AN2 AND2_2407(g17469,g4076,g13217);
  AN2 AND2_2408(g13737,g4501,g10571);
  AN2 AND2_2409(g22038,g5945,g19147);
  AN2 AND2_2410(g23551,g10793,g18948);
  AN2 AND2_2411(g23572,g20230,g20656);
  AN2 AND2_2412(g10917,g9174,g1087);
  AN2 AND2_2413(g12219,g1189,g7532);
  AN2 AND2_2414(g27218,g25997,g16740);
  AN2 AND2_2415(g30927,g29910,g24795);
  AN2 AND2_2416(g18495,g2533,g15426);
  AN2 AND2_2417(g33840,g33253,g20267);
  AN2 AND2_2418(g29641,g28520,g14237);
  AN2 AND2_2419(g29797,g28347,g23259);
  AN2 AND2_2420(g16662,g4552,g14753);
  AN2 AND2_2421(g13697,g11166,g8608);
  AN2 AND2_2422(g28660,g27824,g20623);
  AN2 AND2_2423(g18816,g6527,g15483);
  AN2 AND2_2424(g32011,g8287,g31134);
  AN2 AND2_2425(g27160,g14163,g26340);
  AN2 AND2_2426(g10706,g3338,g8691);
  AN2 AND2_2427(g15113,g4291,g14454);
  AN2 AND2_2428(g19207,g7803,g15992);
  AN2 AND2_2429(g18687,g4664,g15885);
  AN2 AND2_2430(g28456,g27290,g20104);
  AN4 AND4_159(I31097,g32596,g32597,g32598,g32599);
  AN2 AND2_2431(g17601,g9616,g14572);
  AN2 AND2_2432(g22143,g19568,g10971);
  AN2 AND2_2433(g21784,g3423,g20391);
  AN2 AND2_2434(g22937,g753,g20540);
  AN2 AND2_2435(g26845,g24391,g21426);
  AN2 AND2_2436(g14256,g2079,g11872);
  AN2 AND2_2437(g21956,g5360,g21514);
  AN2 AND2_2438(g18752,g15146,g17926);
  AN2 AND2_2439(g27455,g26488,g17603);
  AN2 AND2_2440(g26395,g22547,g25561);
  AN2 AND2_2441(g30604,g18911,g29878);
  AN3 AND3_153(g33522,g32902,I31306,I31307);
  AN2 AND2_2442(g18374,g1878,g15171);
  AN2 AND2_2443(g29635,g28910,g22432);
  AN2 AND2_2444(g21889,g4169,g19801);
  AN2 AND2_2445(g23103,g10143,g20765);
  AN4 AND4_160(g27617,g23032,g26264,g26424,g24982);
  AN2 AND2_2446(g15105,g4235,g14454);
  AN2 AND2_2447(g21980,g5567,g19074);
  AN2 AND2_2448(g10624,g8387,g3072);
  AN2 AND2_2449(g28550,g12009,g27092);
  AN2 AND2_2450(g18643,g3849,g17096);
  AN2 AND2_2451(g7469,g4382,g4438);
  AN2 AND2_2452(g32310,g27577,g31376);
  AN2 AND2_2453(g16204,g6537,g14348);
  AN2 AND2_2454(g28314,g27552,g14205);
  AN2 AND2_2455(g21888,g4165,g19801);
  AN2 AND2_2456(g21824,g3706,g20453);
  AN2 AND2_2457(g26633,g24964,g20616);
  AN2 AND2_2458(g34563,g34372,g17465);
  AN3 AND3_154(I17542,g13156,g6767,g6756);
  AN2 AND2_2459(g27201,g25997,g16685);
  AN2 AND2_2460(g27277,g26359,g14191);
  AN4 AND4_161(I24675,g24022,g24023,g24024,g24025);
  AN3 AND3_155(g33483,g32621,I31111,I31112);
  AN2 AND2_2461(g26719,g10709,g24438);
  AN2 AND2_2462(g24289,g4427,g22550);
  AN2 AND2_2463(g18669,g4608,g17367);
  AN2 AND2_2464(g32112,g31646,g29923);
  AN2 AND2_2465(g25927,g25004,g20375);
  AN2 AND2_2466(g32050,g11003,g30825);
  AN2 AND2_2467(g24309,g4480,g22228);
  AN2 AND2_2468(g33862,g33272,g20504);
  AN2 AND2_2469(g18260,g1252,g16000);
  AN2 AND2_2470(g28243,g27879,g23423);
  AN2 AND2_2471(g24288,g4417,g22550);
  AN2 AND2_2472(g27595,g26733,g26703);
  AN2 AND2_2473(g24224,g269,g22594);
  AN2 AND2_2474(g18668,g4322,g17367);
  AN2 AND2_2475(g27467,g269,g26832);
  AN4 AND4_162(g27494,g8038,g26314,g518,g9077);
  AN2 AND2_2476(g31949,g1287,g30825);
  AN2 AND2_2477(g18392,g1988,g15171);
  AN2 AND2_2478(g29891,g28420,g23356);
  AN2 AND2_2479(g24308,g4489,g22228);
  AN2 AND2_2480(g21931,g5188,g18997);
  AN2 AND2_2481(g18195,g847,g17821);
  AN2 AND2_2482(g22015,g5719,g21562);
  AN2 AND2_2483(g18489,g2509,g15426);
  AN2 AND2_2484(g34395,g34193,g21336);
  AN2 AND2_2485(g31948,g30670,g18884);
  AN2 AND2_2486(g32096,g31601,g29893);
  AN2 AND2_2487(g28269,g27205,g19712);
  AN2 AND2_2488(g29575,g2066,g28604);
  AN2 AND2_2489(g15881,g3582,g13983);
  AN2 AND2_2490(g18559,g12856,g15277);
  AN2 AND2_2491(g25491,g23615,g21355);
  AN2 AND2_2492(g18525,g2610,g15509);
  AN2 AND2_2493(g18488,g2495,g15426);
  AN2 AND2_2494(g18424,g2165,g18008);
  AN2 AND2_2495(g28341,g27240,g19790);
  AN2 AND2_2496(g29711,g2541,g29134);
  AN2 AND2_2497(g33904,g33321,g21059);
  AN2 AND2_2498(g24495,g6928,g23127);
  AN2 AND2_2499(g28268,g8572,g27990);
  AN2 AND2_2500(g31252,g29643,g20101);
  AN2 AND2_2501(g29327,g29070,g22156);
  AN2 AND2_2502(g26861,g25021,g25003);
  AN2 AND2_2503(g33252,g32155,g20064);
  AN2 AND2_2504(g13080,g6923,g11357);
  AN2 AND2_2505(g18558,g2803,g15277);
  AN2 AND2_2506(g28655,g27561,g20603);
  AN2 AND2_2507(g30191,g28647,g23843);
  AN2 AND2_2508(g16233,g6137,g14251);
  AN2 AND2_2509(g29537,g28976,g22472);
  AN2 AND2_2510(g34191,g33713,g24404);
  AN2 AND2_2511(g16672,g6295,g15008);
  AN2 AND2_2512(g27822,g4157,g25893);
  AN4 AND4_163(I27539,g28040,g24135,g24136,g24137);
  AN2 AND2_2513(g26389,g19949,g25553);
  AN2 AND2_2514(g18893,g16215,g16030);
  AN2 AND2_2515(g25981,g2051,g25007);
  AN2 AND2_2516(g24687,g5827,g23666);
  AN4 AND4_164(I31011,g30735,g31797,g32471,g32472);
  AN2 AND2_2517(g27266,g26789,g26770);
  AN2 AND2_2518(g26612,g901,g24407);
  AN4 AND4_165(I27538,g21209,g24132,g24133,g24134);
  AN2 AND2_2519(g26388,g19595,g25552);
  AN2 AND2_2520(g18544,g2791,g15277);
  AN2 AND2_2521(g26324,g2661,g25439);
  AN2 AND2_2522(g32428,g31133,g16261);
  AN2 AND2_2523(g29606,g28480,g8011);
  AN2 AND2_2524(g21024,g16306,g4871);
  AN2 AND2_2525(g18713,g4836,g15915);
  AN2 AND2_2526(g13461,g2719,g11819);
  AN2 AND2_2527(g22084,g6291,g19210);
  AN2 AND2_2528(g31183,g30249,g25174);
  AN2 AND2_2529(g26251,g1988,g25341);
  AN2 AND2_2530(g22110,g15167,g19277);
  AN2 AND2_2531(g24643,g22636,g19696);
  AN2 AND2_2532(g26272,g2036,g25470);
  AN2 AND2_2533(g33847,g33260,g20383);
  AN2 AND2_2534(g21860,g3945,g21070);
  AN2 AND2_2535(g16513,g8345,g13708);
  AN2 AND2_2536(g28694,g27579,g20664);
  AN2 AND2_2537(g29750,g28296,g23215);
  AN2 AND2_2538(g29982,g23656,g28998);
  AN2 AND2_2539(g29381,g28135,g19399);
  AN2 AND2_2540(g18610,g15088,g17059);
  AN2 AND2_2541(g34861,g16540,g34827);
  AN2 AND2_2542(g30247,g28735,g23937);
  AN2 AND2_2543(g18705,g4801,g16782);
  AN2 AND2_2544(g13887,g5204,g12402);
  AN2 AND2_2545(g25990,g9461,g25017);
  AN2 AND2_2546(g23497,g20169,g20569);
  AN3 AND3_156(g33509,g32809,I31241,I31242);
  AN2 AND2_2547(g24669,g22653,g19742);
  AN2 AND2_2548(g31933,g939,g30735);
  AN2 AND2_2549(g30926,g29903,g21163);
  AN2 AND2_2550(g30045,g29200,g12419);
  AN2 AND2_2551(g18255,g1087,g16897);
  AN2 AND2_2552(g18189,g812,g17821);
  AN2 AND2_2553(g27588,g26690,g26673);
  AN2 AND2_2554(g15779,g13909,g11214);
  AN2 AND2_2555(g18679,g4633,g15758);
  AN2 AND2_2556(g31508,g29813,g23459);
  AN2 AND2_2557(g34389,g34170,g20715);
  AN2 AND2_2558(g17321,g1418,g13105);
  AN4 AND4_166(I31112,g32617,g32618,g32619,g32620);
  AN2 AND2_2559(g34045,g33766,g22942);
  AN2 AND2_2560(g30612,g26338,g29597);
  AN3 AND3_157(g33508,g32802,I31236,I31237);
  AN2 AND2_2561(g24668,g11754,g22979);
  AN2 AND2_2562(g21700,g150,g20283);
  AN2 AND2_2563(g30099,g28549,g20776);
  AN2 AND2_2564(g33872,g33282,g20548);
  AN2 AND2_2565(g18270,g1291,g16031);
  AN2 AND2_2566(g29796,g28345,g23258);
  AN2 AND2_2567(g17179,g1041,g13211);
  AN2 AND2_2568(g24392,g3115,g23067);
  AN2 AND2_2569(g22685,g11891,g20192);
  AN2 AND2_2570(g18188,g807,g17328);
  AN2 AND2_2571(g18124,g102,g16886);
  AN2 AND2_2572(g21987,g5579,g19074);
  AN2 AND2_2573(g18678,g66,g15758);
  AN2 AND2_2574(g34388,g10802,g34062);
  AN2 AND2_2575(g16026,g854,g14065);
  AN2 AND2_2576(g28557,g27772,g15647);
  AN2 AND2_2577(g34324,g14064,g34161);
  AN2 AND2_2578(g15081,g2689,g12983);
  AN2 AND2_2579(g13393,g703,g11048);
  AN2 AND2_2580(g16212,g6167,g14321);
  AN2 AND2_2581(g24195,g74,g22722);
  AN2 AND2_2582(g28210,g9229,g27554);
  AN2 AND2_2583(g32317,g5507,g31542);
  AN2 AND2_2584(g27119,g25877,g22542);
  AN2 AND2_2585(g30098,g28548,g20774);
  AN2 AND2_2586(g34701,g34536,g20179);
  AN4 AND4_167(g10721,g3288,g6875,g3274,g8481);
  AN2 AND2_2587(g20559,g336,g15831);
  AN2 AND2_2588(g30251,g28745,g23940);
  AN2 AND2_2589(g34534,g34321,g19743);
  AN2 AND2_2590(g23658,g14687,g20852);
  AN2 AND2_2591(g30272,g28814,g23982);
  AN3 AND3_158(g34098,g33744,g9104,g18957);
  AN2 AND2_2592(g19206,g460,g16206);
  AN2 AND2_2593(g15786,g13940,g11233);
  AN2 AND2_2594(g18460,g2351,g15224);
  AN2 AND2_2595(g18686,g4659,g15885);
  AN2 AND2_2596(g24559,g22993,g19567);
  AN2 AND2_2597(g18383,g1950,g15171);
  AN2 AND2_2598(g29840,g2153,g29056);
  AN2 AND2_2599(g24488,g6905,g23082);
  AN4 AND4_168(I31096,g31376,g31812,g32594,g32595);
  AN2 AND2_2600(g24016,g14528,g21610);
  AN2 AND2_2601(g27118,g26055,g16529);
  AN3 AND3_159(g22417,g7753,g9285,g21186);
  AN2 AND2_2602(g11960,g2495,g7424);
  AN2 AND2_2603(g32129,g31658,g29955);
  AN2 AND2_2604(g21943,g5240,g18997);
  AN2 AND2_2605(g25832,g8219,g24625);
  AN2 AND2_2606(g21296,g7879,g16072);
  AN2 AND2_2607(g24558,g22516,g19566);
  AN2 AND2_2608(g18267,g1266,g16000);
  AN2 AND2_2609(g18294,g15072,g16449);
  AN2 AND2_2610(g27616,g26349,g20449);
  AN2 AND2_2611(g26871,g25038,g25020);
  AN2 AND2_2612(g17654,g962,g13284);
  AN2 AND2_2613(g32128,g31631,g29953);
  AN3 AND3_160(I17575,g13156,g11450,g6756);
  AN2 AND2_2614(g27313,g1982,g26701);
  AN2 AND2_2615(g29192,g27163,g10290);
  AN2 AND2_2616(g30032,g29072,g9326);
  AN2 AND2_2617(g21969,g5373,g21514);
  AN2 AND2_2618(g26360,g10589,g25533);
  AN2 AND2_2619(g25573,I24704,I24705);
  AN2 AND2_2620(g30140,g28600,g23749);
  AN2 AND2_2621(g27276,g9750,g26607);
  AN2 AND2_2622(g27285,g9912,g26632);
  AN2 AND2_2623(g29522,g28923,g22369);
  AN2 AND2_2624(g32323,g31311,g20610);
  AN2 AND2_2625(g24865,g11323,g23253);
  AN2 AND2_2626(g29663,g1950,g28693);
  AN2 AND2_2627(g34140,g33931,g23802);
  AN2 AND2_2628(g22762,g9305,g20645);
  AN2 AND2_2629(g15651,g429,g13414);
  AN2 AND2_2630(g21968,g5459,g21514);
  AN2 AND2_2631(g10655,g8440,g3423);
  AN2 AND2_2632(g15672,g433,g13458);
  AN2 AND2_2633(g27305,g10041,g26683);
  AN2 AND2_2634(g25926,g25005,g24839);
  AN2 AND2_2635(g24713,g5831,g23666);
  AN2 AND2_2636(g25045,g17525,g23448);
  AN2 AND2_2637(g18219,g969,g16100);
  AN2 AND2_2638(g27254,g25935,g19688);
  AN2 AND2_2639(g30061,g1036,g28188);
  AN2 AND2_2640(g33311,g31942,g12925);
  AN2 AND2_2641(g21855,g3925,g21070);
  AN2 AND2_2642(g34061,g33800,g23076);
  AN2 AND2_2643(g14180,g872,g10632);
  AN2 AND2_2644(g23855,g4112,g19455);
  AN2 AND2_2645(g22216,g13660,g20000);
  AN2 AND2_2646(g18218,g1008,g16100);
  AN2 AND2_2647(g21870,g4093,g19801);
  AN3 AND3_161(I17606,g14988,g11450,g6756);
  AN2 AND2_2648(g28601,g27506,g20514);
  AN2 AND2_2649(g28677,g27571,g20635);
  AN2 AND2_2650(g27036,g26329,g11038);
  AN2 AND2_2651(g29553,g2437,g28911);
  AN2 AND2_2652(g26629,g14173,g24418);
  AN2 AND2_2653(g27177,g25997,g16651);
  AN2 AND2_2654(g27560,g26299,g20191);
  AN2 AND2_2655(g34871,g34823,g19908);
  AN2 AND2_2656(g24189,g324,g22722);
  AN2 AND2_2657(g31756,g30114,g23942);
  AN2 AND2_2658(g24679,g13289,g22985);
  AN2 AND2_2659(g11244,g8346,g8566);
  AN2 AND2_2660(g29949,g23575,g28924);
  AN2 AND2_2661(g32232,g31241,g20266);
  AN2 AND2_2662(g20188,g5849,g17772);
  AN2 AND2_2663(g18160,g645,g17433);
  AN2 AND2_2664(g29326,g29105,g22155);
  AN3 AND3_162(g10838,g7738,g5527,g5535);
  AN2 AND2_2665(g28143,g27344,g26083);
  AN2 AND2_2666(g31780,g30163,g23999);
  AN3 AND3_163(g25462,g6404,g22300,I24585);
  AN2 AND2_2667(g24188,g316,g22722);
  AN2 AND2_2668(g22117,g6597,g19277);
  AN2 AND2_2669(g29536,g28969,g22432);
  AN2 AND2_2670(g22000,g5727,g21562);
  AN2 AND2_2671(g21867,g4082,g19801);
  AN2 AND2_2672(g18455,g2327,g15224);
  AN2 AND2_2673(g24686,g5485,g23630);
  AN2 AND2_2674(g24939,g23771,g21012);
  AN2 AND2_2675(g29757,g28305,g23221);
  AN4 AND4_169(I31317,g32914,g32915,g32916,g32917);
  AN2 AND2_2676(g33350,g32235,g20702);
  AN2 AND2_2677(g32261,g31251,g20386);
  AN2 AND2_2678(g18617,g3462,g17062);
  AN2 AND2_2679(g18470,g2403,g15224);
  AN2 AND2_2680(g20093,g15372,g14584);
  AN2 AND2_2681(g33820,g33075,g26830);
  AN2 AND2_2682(g29621,g2449,g28994);
  AN3 AND3_164(I24576,g5390,g5396,g9792);
  AN3 AND3_165(I24585,g9621,g9892,g6439);
  AN2 AND2_2683(g10619,g3080,g7907);
  AN2 AND2_2684(g21714,g278,g20283);
  AN2 AND2_2685(g23581,g20183,g11900);
  AN2 AND2_2686(g24294,g4452,g22550);
  AN2 AND2_2687(g31152,g10039,g30067);
  AN2 AND2_2688(g25061,g17586,g23461);
  AN4 AND4_170(I31002,g32459,g32460,g32461,g32462);
  AN2 AND2_2689(g18201,g15061,g15938);
  AN2 AND2_2690(g33846,g33259,g20380);
  AN4 AND4_171(I31057,g32538,g32539,g32540,g32541);
  AN2 AND2_2691(g21707,g191,g20283);
  AN2 AND2_2692(g21819,g3614,g20924);
  AN2 AND2_2693(g29564,g1882,g28896);
  AN2 AND2_2694(g18277,g1312,g16136);
  AN2 AND2_2695(g14210,g4392,g10590);
  AN2 AND2_2696(g21910,g5016,g21468);
  AN2 AND2_2697(g26147,g6513,g25133);
  AN2 AND2_2698(g30220,g28699,g23888);
  AN2 AND2_2699(g28666,g27567,g20625);
  AN2 AND2_2700(g33731,g33116,g19520);
  AN2 AND2_2701(g28217,g27733,g23391);
  AN2 AND2_2702(g22123,g6609,g19277);
  AN2 AND2_2703(g21818,g3610,g20924);
  AN4 AND4_172(g17747,g6772,g11592,g11640,I18740);
  AN2 AND2_2704(g21979,g5559,g19074);
  AN2 AND2_2705(g16896,g262,g13120);
  AN2 AND2_2706(g27665,g26872,g23519);
  AN2 AND2_2707(g30246,g28734,g23936);
  AN2 AND2_2708(g25871,g8334,g24804);
  AN2 AND2_2709(g20875,g16281,g4681);
  AN2 AND2_2710(g18595,g2927,g16349);
  AN2 AND2_2711(g28478,g27007,g12345);
  AN2 AND2_2712(g18467,g2380,g15224);
  AN2 AND2_2713(g18494,g2527,g15426);
  AN2 AND2_2714(g19500,g504,g16712);
  AN2 AND2_2715(g24219,g225,g22594);
  AN2 AND2_2716(g26858,g2970,g24540);
  AN2 AND2_2717(g21978,g5551,g19074);
  AN2 AND2_2718(g11967,g311,g7802);
  AN2 AND2_2719(g18623,g3484,g17062);
  AN2 AND2_2720(g20218,g6541,g17815);
  AN2 AND2_2721(g30071,g29184,g12975);
  AN2 AND2_2722(g17123,g225,g13209);
  AN2 AND2_2723(g24218,g872,g22594);
  AN2 AND2_2724(g21986,g5575,g19074);
  AN2 AND2_2725(g34071,g8854,g33799);
  AN2 AND2_2726(g18782,g5835,g18065);
  AN2 AND2_2727(g27485,g26519,g17644);
  AN2 AND2_2728(g28556,g27431,g20374);
  AN2 AND2_2729(g29509,g1600,g28755);
  AN2 AND2_2730(g32316,g31307,g23522);
  AN2 AND2_2731(g33405,g32354,g21398);
  AN2 AND2_2732(g21741,g15086,g20330);
  AN2 AND2_2733(g26844,g25261,g21418);
  AN2 AND2_2734(g18419,g2051,g15373);
  AN2 AND2_2735(g27454,g26488,g17602);
  AN2 AND2_2736(g26394,g22530,g25560);
  AN2 AND2_2737(g18352,g1798,g17955);
  AN2 AND2_2738(g29634,g2108,g29121);
  AN2 AND2_2739(g29851,g1668,g29079);
  AN2 AND2_2740(g29872,g28401,g23333);
  AN2 AND2_2741(g28223,g27338,g17194);
  AN2 AND2_2742(g15104,g6955,g14454);
  AN2 AND2_2743(g34754,g34677,g19602);
  AN2 AND2_2744(g18155,g15056,g17533);
  AN2 AND2_2745(g21067,g10085,g17625);
  AN2 AND2_2746(g18418,g2122,g15373);
  AN2 AND2_2747(g18822,g6723,g15680);
  AN2 AND2_2748(g30825,g29814,g22332);
  AN2 AND2_2749(g19613,g1437,g16713);
  AN2 AND2_2750(g32056,g27271,g31021);
  AN2 AND2_2751(g18266,g1274,g16000);
  AN2 AND2_2752(g11010,g4698,g8933);
  AN2 AND2_2753(g34859,g16540,g34820);
  AN2 AND2_2754(g18170,g661,g17433);
  AN4 AND4_173(I31232,g32791,g32792,g32793,g32794);
  AN2 AND2_2755(g10677,g4141,g7611);
  AN2 AND2_2756(g22992,g1227,g19765);
  AN2 AND2_2757(g34370,g34067,g10554);
  AN4 AND4_174(I24674,g19919,g24019,g24020,g24021);
  AN2 AND2_2758(g21801,g3554,g20924);
  AN2 AND2_2759(g28110,g27974,g18886);
  AN2 AND2_2760(g21735,g3057,g20330);
  AN2 AND2_2761(g21877,g6888,g19801);
  AN2 AND2_2762(g23801,g1448,g19362);
  AN2 AND2_2763(g34858,g16540,g34816);
  AN2 AND2_2764(g30151,g28607,g21249);
  AN2 AND2_2765(g30172,g28625,g21286);
  AN2 AND2_2766(g24915,g23087,g20158);
  AN4 AND4_175(I31261,g30937,g31842,g32831,g32832);
  AN2 AND2_2767(g27594,g26721,g26694);
  AN2 AND2_2768(g28531,g27722,g15608);
  AN2 AND2_2769(g17391,g9556,g14378);
  AN2 AND2_2770(g22835,g15803,g19633);
  AN2 AND2_2771(g28178,g27019,g19397);
  AN2 AND2_2772(g18167,g718,g17433);
  AN2 AND2_2773(g18194,g843,g17821);
  AN2 AND2_2774(g18589,g2902,g16349);
  AN2 AND2_2775(g22014,g5805,g21562);
  AN2 AND2_2776(g34367,g7404,g34042);
  AN2 AND2_2777(g31787,g21281,g29385);
  AN2 AND2_2778(g34394,g34190,g21305);
  AN2 AND2_2779(g25071,g12804,g23478);
  AN2 AND2_2780(g33113,g31964,g22339);
  AN2 AND2_2781(g33787,g33103,g20595);
  AN2 AND2_2782(g32342,g6545,g31579);
  AN2 AND2_2783(g29574,g2016,g28931);
  AN2 AND2_2784(g31282,g30130,g27779);
  AN2 AND2_2785(g22007,g5770,g21562);
  AN2 AND2_2786(g15850,g3606,g14151);
  AN3 AND3_166(g29205,g24117,I27523,I27524);
  AN2 AND2_2787(g18588,g2970,g16349);
  AN2 AND2_2788(g18524,g2681,g15509);
  AN2 AND2_2789(g28676,g27570,g20632);
  AN2 AND2_2790(g32145,g31609,g29977);
  AN2 AND2_2791(g14791,g1146,g10909);
  AN2 AND2_2792(g32031,g31372,g13464);
  AN2 AND2_2793(g24467,g13761,g23047);
  AN2 AND2_2794(g27519,g26488,g17710);
  AN2 AND2_2795(g33357,g32247,g20775);
  AN3 AND3_167(g27185,g26190,g8302,g1917);
  AN2 AND2_2796(g25147,g20202,g23542);
  AN2 AND2_2797(g32199,g30916,g25506);
  AN2 AND2_2798(g18401,g2036,g15373);
  AN2 AND2_2799(g28654,g1030,g27108);
  AN2 AND2_2800(g33105,g26298,g32138);
  AN2 AND2_2801(g14168,g887,g10632);
  AN2 AND2_2802(g18477,g2429,g15426);
  AN2 AND2_2803(g26203,g1632,g25337);
  AN2 AND2_2804(g33743,g33119,g19574);
  AN2 AND2_2805(g16802,g5567,g14807);
  AN2 AND2_2806(g18119,g475,g17015);
  AN2 AND2_2807(g27518,g26488,g17709);
  AN2 AND2_2808(g27154,g26055,g16630);
  AN2 AND2_2809(g34319,g9535,g34156);
  AN2 AND2_2810(g32198,g4253,g31327);
  AN2 AND2_2811(g22116,g6589,g19277);
  AN2 AND2_2812(g16730,g5212,g14723);
  AN2 AND2_2813(g24984,g22929,g12818);
  AN2 AND2_2814(g18118,g471,g17015);
  AN2 AND2_2815(g21866,g4072,g19801);
  AN2 AND2_2816(g21917,g5092,g21468);
  AN2 AND2_2817(g30227,g28708,g23899);
  AN2 AND2_2818(g31769,g30141,g23986);
  AN2 AND2_2819(g23917,g1472,g19428);
  AN2 AND2_2820(g33640,g33387,g18831);
  AN4 AND4_176(g26281,g24688,g8812,g8778,g8757);
  AN2 AND2_2821(g32330,g31320,g20631);
  AN2 AND2_2822(g29592,g28469,g11832);
  AN2 AND2_2823(g30059,g28106,g12467);
  AN2 AND2_2824(g22720,g9253,g20619);
  AN4 AND4_177(I31316,g29385,g32911,g32912,g32913);
  AN2 AND2_2825(g30025,g28492,g23502);
  AN2 AND2_2826(g25151,g17719,g23549);
  AN2 AND2_2827(g16765,g6581,g15045);
  AN2 AND2_2828(g15716,g468,g13437);
  AN2 AND2_2829(g18749,g5148,g17847);
  AN2 AND2_2830(g22041,g5957,g19147);
  AN2 AND2_2831(g26301,g2145,g25244);
  AN2 AND2_2832(g13656,g278,g11144);
  AN2 AND2_2833(g18616,g6875,g17200);
  AN2 AND2_2834(g18313,g1430,g16931);
  AN2 AND2_2835(g33803,g33231,g20071);
  AN3 AND3_168(g24822,g3010,g23534,I24003);
  AN2 AND2_2836(g26120,g9809,g25293);
  AN2 AND2_2837(g30058,g29180,g12950);
  AN2 AND2_2838(g16690,g8399,g13867);
  AN4 AND4_178(g11144,g239,g8136,g246,I14198);
  AN2 AND2_2839(g18748,g5142,g17847);
  AN2 AND2_2840(g8643,g2927,g2922);
  AN2 AND2_2841(g25367,g6946,g22407);
  AN4 AND4_179(I31056,g30735,g31805,g32536,g32537);
  AN2 AND2_2842(g21706,g222,g20283);
  AN2 AND2_2843(g18276,g1351,g16136);
  AN2 AND2_2844(g18285,g1395,g16164);
  AN2 AND2_2845(g29350,g4939,g28395);
  AN2 AND2_2846(g26146,g9892,g25334);
  AN2 AND2_2847(g30203,g28668,g23864);
  AN2 AND2_2848(g18704,g4793,g16782);
  AN2 AND2_2849(g34203,g33726,g24537);
  AN2 AND2_2850(g18305,g1521,g16489);
  AN2 AND2_2851(g33881,g33292,g20586);
  AN2 AND2_2852(g30044,g29174,g12944);
  AN2 AND2_2853(g18254,g1236,g16897);
  AN2 AND2_2854(g18809,g7074,g15656);
  AN2 AND2_2855(g21923,g5029,g21468);
  AN2 AND2_2856(g22340,g19605,g13522);
  AN2 AND2_2857(g32161,g3151,g31154);
  AN2 AND2_2858(g22035,g5933,g19147);
  AN2 AND2_2859(g28587,g27487,g20498);
  AN2 AND2_2860(g26290,g2595,g25498);
  AN2 AND2_2861(g18466,g2389,g15224);
  AN2 AND2_2862(g23280,g19417,g20146);
  AN2 AND2_2863(g27215,g26055,g16724);
  AN2 AND2_2864(g27501,g26400,g17673);
  AN2 AND2_2865(g15112,g4284,g14454);
  AN4 AND4_180(I31271,g29385,g32846,g32847,g32848);
  AN2 AND2_2866(g30281,g28850,g23992);
  AN2 AND2_2867(g18808,g6390,g15656);
  AN3 AND3_169(g25420,g6058,g22220,I24555);
  AN2 AND2_2868(g24194,g106,g22722);
  AN2 AND2_2869(g24589,g5471,g23630);
  AN2 AND2_2870(g34281,g34043,g19276);
  AN2 AND2_2871(g29731,g2089,g29118);
  AN2 AND2_2872(g22142,g7957,g19140);
  AN2 AND2_2873(g27439,g232,g26831);
  AN2 AND2_2874(g34301,g34064,g19415);
  AN2 AND2_2875(g18177,g749,g17328);
  AN2 AND2_2876(g18560,g2837,g15277);
  AN2 AND2_2877(g30120,g28576,g21051);
  AN2 AND2_2878(g28543,g27735,g15628);
  AN2 AND2_2879(g24588,g5142,g23590);
  AN2 AND2_2880(g32087,g1291,g30825);
  AN2 AND2_2881(g34120,g33930,g25158);
  AN4 AND4_181(I31342,g32949,g32950,g32951,g32952);
  AN2 AND2_2882(g32258,g31624,g30303);
  AN2 AND2_2883(g28117,g8075,g27245);
  AN2 AND2_2884(g18642,g15097,g17096);
  AN2 AND2_2885(g25059,g20870,g23460);
  AN2 AND2_2886(g33890,g33310,g20659);
  AN2 AND2_2887(g19788,g9983,g17216);
  AN4 AND4_182(I31031,g30614,g31801,g32499,g32500);
  AN2 AND2_2888(g16128,g14333,g14166);
  AN2 AND2_2889(g34146,g33788,g20091);
  AN2 AND2_2890(g34738,g34660,g33442);
  AN2 AND2_2891(g33249,g32144,g20026);
  AN2 AND2_2892(g34562,g34369,g17411);
  AN2 AND2_2893(g28569,g27453,g20433);
  AN2 AND2_2894(g21066,g10043,g17625);
  AN2 AND2_2895(g25058,g23276,g20513);
  AN2 AND2_2896(g16245,g14278,g14708);
  AN2 AND2_2897(g32043,g31482,g16173);
  AN3 AND3_170(g33482,g32614,I31106,I31107);
  AN2 AND2_2898(g32244,g31609,g30297);
  AN2 AND2_2899(g31710,g29814,g19128);
  AN2 AND2_2900(g33248,g32131,g19996);
  AN2 AND2_2901(g10676,g8506,g3774);
  AN4 AND4_183(I27514,g24091,g24092,g24093,g24094);
  AN2 AND2_2902(g18733,g15141,g16877);
  AN2 AND2_2903(g27083,g25819,g22456);
  AN2 AND2_2904(g27348,g26488,g17392);
  AN2 AND2_2905(g33710,g14037,g33246);
  AN2 AND2_2906(g22130,g6637,g19277);
  AN2 AND2_2907(g27284,g9908,g26631);
  AN2 AND2_2908(g24864,g11201,g22305);
  AN2 AND2_2909(g22193,g19880,g20682);
  AN2 AND2_2910(g28242,g27769,g23626);
  AN2 AND2_2911(g21876,g4119,g19801);
  AN2 AND2_2912(g21885,g4122,g19801);
  AN2 AND2_2913(g26547,g13283,g25027);
  AN2 AND2_2914(g10654,g3085,g8434);
  AN2 AND2_2915(g11023,g9669,g5084);
  AN2 AND2_2916(g15857,g3199,g14038);
  AN2 AND2_2917(g23885,g4132,g19513);
  AN2 AND2_2918(g27304,g2273,g26682);
  AN2 AND2_2919(g24749,g17511,g22432);
  AN2 AND2_2920(g32069,g10878,g30735);
  AN2 AND2_2921(g12284,g1532,g7557);
  AN2 AND2_2922(g14654,g7178,g10476);
  AN2 AND2_2923(g24313,g4504,g22228);
  AN2 AND2_2924(g22165,g15594,g18903);
  AN2 AND2_2925(g18630,g3689,g17226);
  AN2 AND2_2926(g21854,g3921,g21070);
  AN2 AND2_2927(g15793,g3219,g13873);
  AN2 AND2_2928(g18693,g4717,g16053);
  AN2 AND2_2929(g23854,g4093,g19506);
  AN2 AND2_2930(g31778,g21369,g29385);
  AN2 AND2_2931(g24748,g17656,g22457);
  AN4 AND4_184(g26226,g24688,g8812,g10658,g10627);
  AN2 AND2_2932(g32068,g31515,g10862);
  AN2 AND2_2933(g33081,g32388,g18875);
  AN2 AND2_2934(g17193,g2504,g13023);
  AN2 AND2_2935(g21763,g3223,g20785);
  AN2 AND2_2936(g18166,g655,g17433);
  AN2 AND2_2937(g24285,g4388,g22550);
  AN2 AND2_2938(g25902,g24398,g19373);
  AN2 AND2_2939(g18665,g4584,g17367);
  AN4 AND4_185(I31132,g32645,g32646,g32647,g32648);
  AN2 AND2_2940(g31786,g30189,g24010);
  AN2 AND2_2941(g25957,g17190,g24960);
  AN2 AND2_2942(g24704,g17593,g22384);
  AN3 AND3_171(g25377,g5712,g22210,I24530);
  AN2 AND2_2943(g33786,g33130,g20572);
  AN2 AND2_2944(g24305,g4477,g22228);
  AN2 AND2_2945(g16737,g6645,g15042);
  AN2 AND2_2946(g26572,g7443,g24439);
  AN2 AND2_2947(g22006,g5767,g21562);
  AN2 AND2_2948(g28639,g27767,g20597);
  AN3 AND3_172(g24900,g3752,g23582,I24067);
  AN2 AND2_2949(g33647,g33390,g18878);
  AN2 AND2_2950(g32337,g31465,g20663);
  AN2 AND2_2951(g27139,g26055,g16608);
  AN3 AND3_173(g28293,g7424,g2495,g27474);
  AN2 AND2_2952(g33356,g32245,g20772);
  AN2 AND2_2953(g22863,g9547,g20388);
  AN2 AND2_2954(g27653,g26549,g15562);
  AN2 AND2_2955(g28638,g27551,g20583);
  AN2 AND2_2956(g32171,g31706,g27800);
  AN4 AND4_186(I31161,g30614,g31824,g32687,g32688);
  AN2 AND2_2957(g18476,g2433,g15426);
  AN2 AND2_2958(g18485,g2465,g15426);
  AN2 AND2_2959(g29787,g28334,g23249);
  AN2 AND2_2960(g26127,g2236,g25119);
  AN2 AND2_2961(g27138,g26055,g16607);
  AN2 AND2_2962(g28265,g11367,g27989);
  AN2 AND2_2963(g34661,g34575,g18907);
  AN2 AND2_2964(g18555,g2834,g15277);
  AN2 AND2_2965(g18454,g2303,g15224);
  AN3 AND3_174(g25290,g5022,g22173,I24482);
  AN2 AND2_2966(g14216,g7631,g10608);
  AN2 AND2_2967(g21916,g5084,g21468);
  AN2 AND2_2968(g30226,g28707,g23898);
  AN2 AND2_2969(g18570,g2848,g16349);
  AN2 AND2_2970(g18712,g4843,g15915);
  AN2 AND2_2971(g33233,g32094,g23005);
  AN2 AND2_2972(g31182,g30240,g20682);
  AN2 AND2_2973(g31672,g29814,g19050);
  AN2 AND2_2974(g27333,g10180,g26765);
  AN2 AND2_2975(g24642,g8290,g22898);
  AN2 AND2_2976(g34226,g33914,g21467);
  AN2 AND2_2977(g14587,g10584,g10567);
  AN2 AND2_2978(g29743,g28206,g10233);
  AN4 AND4_187(I31087,g32580,g32581,g32582,g32583);
  AN2 AND2_2979(g34715,g34570,g33375);
  AN2 AND2_2980(g34481,g34404,g18916);
  AN2 AND2_2981(g23314,g9104,g19200);
  AN2 AND2_2982(g32425,g31668,g21604);
  AN2 AND2_2983(g26103,g2185,g25100);
  AN2 AND2_2984(g34572,g34387,g33326);
  AN2 AND2_2985(g10543,g8238,g437);
  AN2 AND2_2986(g26095,g11923,g25090);
  AN2 AND2_2987(g27963,g25952,g16047);
  AN2 AND2_2988(g23076,g19128,g9104);
  AN2 AND2_2989(g29640,g28498,g8125);
  AN2 AND2_2990(g25366,g7733,g22406);
  AN2 AND2_2991(g29769,g28319,g23237);
  AN2 AND2_2992(g18239,g1135,g16326);
  AN2 AND2_2993(g21721,g385,g21037);
  AN2 AND2_2994(g33331,g32216,g20607);
  AN2 AND2_2995(g27664,g1024,g25911);
  AN2 AND2_2996(g18567,g2894,g16349);
  AN2 AND2_2997(g18594,g12858,g16349);
  AN2 AND2_2998(g31513,g2606,g29318);
  AN2 AND2_2999(g32010,g31785,g22303);
  AN3 AND3_175(g33513,g32837,I31261,I31262);
  AN2 AND2_3000(g29803,g28414,g26836);
  AN2 AND2_3001(g18238,g1152,g16326);
  AN2 AND2_3002(g26181,g2652,g25157);
  AN2 AND2_3003(g26671,g316,g24429);
  AN2 AND2_3004(g28586,g27484,g20497);
  AN2 AND2_3005(g24630,g23255,g14149);
  AN2 AND2_3006(g31961,g31751,g22154);
  AN2 AND2_3007(g33897,g33315,g20777);
  AN4 AND4_188(g17781,g6772,g11592,g6789,I18785);
  AN2 AND2_3008(g31505,g30195,g24379);
  AN2 AND2_3009(g28442,g27278,g20072);
  AN3 AND3_176(g33505,g32779,I31221,I31222);
  AN2 AND2_3010(g18382,g1936,g15171);
  AN2 AND2_3011(g24009,g19671,g10971);
  AN2 AND2_3012(g33404,g32353,g21397);
  AN2 AND2_3013(g29881,g2040,g29150);
  AN2 AND2_3014(g21773,g3263,g20785);
  AN2 AND2_3015(g18519,g2648,g15509);
  AN2 AND2_3016(g11016,g4888,g8984);
  AN2 AND2_3017(g21942,g5236,g18997);
  AN2 AND2_3018(g13525,g10019,g11911);
  AN2 AND2_3019(g18176,g732,g17328);
  AN2 AND2_3020(g18185,g790,g17328);
  AN2 AND2_3021(g22063,g6109,g21611);
  AN2 AND2_3022(g18675,g4349,g15758);
  AN2 AND2_3023(g34385,g34168,g20642);
  AN2 AND2_3024(g33717,g14092,g33306);
  AN2 AND2_3025(g24008,g7909,g19502);
  AN2 AND2_3026(g32086,g7597,g30735);
  AN2 AND2_3027(g30095,g28545,g20768);
  AN2 AND2_3028(g31212,g20028,g29669);
  AN2 AND2_3029(g28116,g27366,g26183);
  AN2 AND2_3030(g18518,g2657,g15509);
  AN2 AND2_3031(g18154,g622,g17533);
  AN2 AND2_3032(g27312,g12019,g26700);
  AN2 AND2_3033(g24892,g11559,g23264);
  AN4 AND4_189(g26190,g25357,g11724,g7586,g11686);
  AN2 AND2_3034(g24485,g10710,g22319);
  AN2 AND2_3035(g24476,g18879,g22330);
  AN4 AND4_190(I31337,g32942,g32943,g32944,g32945);
  AN2 AND2_3036(g16611,g5583,g14727);
  AN2 AND2_3037(g27115,g26026,g16526);
  AN2 AND2_3038(g11893,g1668,g7268);
  AN4 AND4_191(g13830,g11543,g11424,g11395,I16143);
  AN2 AND2_3039(g22873,g19854,g19683);
  AN2 AND2_3040(g25551,g23822,g21511);
  AN2 AND2_3041(g18637,g3821,g17096);
  AN2 AND2_3042(g25572,I24699,I24700);
  AN4 AND4_192(I31171,g31528,g31826,g32701,g32702);
  AN2 AND2_3043(g30181,g28636,g23821);
  AN2 AND2_3044(g30671,g29319,g22317);
  AN2 AND2_3045(g18935,g4322,g15574);
  AN2 AND2_3046(g32322,g31308,g20605);
  AN2 AND2_3047(g24555,g23184,g21024);
  AN2 AND2_3048(g29662,g1848,g29049);
  AN2 AND2_3049(g9217,g632,g626);
  AN2 AND2_3050(g21734,g3040,g20330);
  AN2 AND2_3051(g32159,g31658,g30040);
  AN2 AND2_3052(g24712,g19592,g23001);
  AN2 AND2_3053(g29890,g28419,g23355);
  AN2 AND2_3054(g24914,g8721,g23301);
  AN2 AND2_3055(g21839,g3763,g20453);
  AN2 AND2_3056(g21930,g5180,g18997);
  AN2 AND2_3057(g25127,g13997,g23524);
  AN2 AND2_3058(g21993,g5603,g19074);
  AN2 AND2_3059(g32158,g31658,g30022);
  AN2 AND2_3060(g22209,g19907,g20751);
  AN2 AND2_3061(g15856,g9056,g14223);
  AN3 AND3_177(g15995,g13314,g1157,g10666);
  AN2 AND2_3062(g33723,g14091,g33299);
  AN2 AND2_3063(g28237,g9492,g27597);
  AN2 AND2_3064(g21838,g3747,g20453);
  AN2 AND2_3065(g22834,g102,g19630);
  AN2 AND2_3066(g15880,g3211,g13980);
  AN2 AND2_3067(g31149,g29508,g23021);
  AN2 AND2_3068(g21965,g15149,g21514);
  AN2 AND2_3069(g26088,g6545,g25080);
  AN2 AND2_3070(g26024,g2619,g25039);
  AN2 AND2_3071(g22208,g19906,g20739);
  AN2 AND2_3072(g29710,g2380,g29094);
  AN3 AND3_178(g28035,g24103,I26530,I26531);
  AN2 AND2_3073(g29552,g2223,g28579);
  AN2 AND2_3074(g33433,g32238,g29694);
  AN2 AND2_3075(g23131,g13919,g19930);
  AN2 AND2_3076(g32295,g27931,g31376);
  AN2 AND2_3077(g10841,g8509,g8567);
  AN3 AND3_179(g29204,g24110,I27518,I27519);
  AN2 AND2_3078(g31148,g2661,g30055);
  AN2 AND2_3079(g30190,g28646,g23842);
  AN2 AND2_3080(g13042,g433,g11048);
  AN2 AND2_3081(g16199,g3614,g14051);
  AN2 AND2_3082(g18215,g943,g15979);
  AN2 AND2_3083(g25103,g4927,g22908);
  AN2 AND2_3084(g27184,g26628,g13756);
  AN2 AND2_3085(g16736,g6303,g15036);
  AN2 AND2_3086(g18501,g12854,g15509);
  AN2 AND2_3087(g18729,g15139,g16821);
  AN2 AND2_3088(g22021,g5869,g19147);
  AN2 AND2_3089(g27674,g26873,g23543);
  AN2 AND2_3090(g25980,g1926,g25006);
  AN2 AND2_3091(g18577,g2988,g16349);
  AN2 AND2_3092(g33104,g26296,g32137);
  AN2 AND2_3093(g25095,g23319,g20556);
  AN2 AND2_3094(g33811,g33439,g17573);
  AN2 AND2_3095(g33646,g33389,g18876);
  AN2 AND2_3096(g19767,g16810,g14203);
  AN2 AND2_3097(g32336,g31596,g11842);
  AN2 AND2_3098(g34520,g34294,g19505);
  AN2 AND2_3099(g23619,g19453,g13045);
  AN2 AND2_3100(g33343,g32227,g20665);
  AN2 AND2_3101(g21557,g12980,g15674);
  AN2 AND2_3102(g18728,g4939,g16821);
  AN2 AND2_3103(g18439,g2250,g18008);
  AN2 AND2_3104(g30089,g28538,g20709);
  AN2 AND2_3105(g24941,g23171,g20190);
  AN2 AND2_3106(g26126,g1959,g25118);
  AN2 AND2_3107(g30211,g28685,g23878);
  AN2 AND2_3108(g11939,g2361,g7380);
  AN2 AND2_3109(g23618,g19388,g11917);
  AN2 AND2_3110(g25181,g23405,g20696);
  AN3 AND3_180(g34089,g22957,g9104,g33744);
  AN2 AND2_3111(g16843,g6251,g14864);
  AN2 AND2_3112(g18438,g2236,g18008);
  AN2 AND2_3113(g34211,g33891,g21349);
  AN2 AND2_3114(g26250,g1902,g25429);
  AN2 AND2_3115(g13383,g4765,g11797);
  AN2 AND2_3116(g24675,g17568,g22342);
  AN2 AND2_3117(g29647,g28934,g22457);
  AN2 AND2_3118(g30024,g28497,g23501);
  AN2 AND2_3119(g33369,g32277,g21060);
  AN3 AND3_181(I24048,g3034,g3040,g8426);
  AN2 AND2_3120(g17726,g1467,g13315);
  AN2 AND2_3121(g16764,g6307,g14776);
  AN3 AND3_182(g34088,g33736,g9104,g18957);
  AN2 AND2_3122(g13030,g429,g11048);
  AN2 AND2_3123(g22073,g6235,g19210);
  AN2 AND2_3124(g18349,g1768,g17955);
  AN2 AND2_3125(g14586,g11953,g11970);
  AN2 AND2_3126(g13294,g1564,g11513);
  AN4 AND4_193(I31086,g31554,g31811,g32578,g32579);
  AN2 AND2_3127(g29380,g28134,g19396);
  AN2 AND2_3128(g33368,g32275,g21057);
  AN2 AND2_3129(g34860,g16540,g34823);
  AN2 AND2_3130(g16869,g6259,g14902);
  AN2 AND2_3131(g27692,g26392,g20697);
  AN2 AND2_3132(g28130,g27353,g23063);
  AN2 AND2_3133(g28193,g8851,g27629);
  AN2 AND2_3134(g26339,g225,g24836);
  AN2 AND2_3135(g25931,g24574,g19477);
  AN2 AND2_3136(g18906,g13568,g16264);
  AN2 AND2_3137(g18348,g1744,g17955);
  AN2 AND2_3138(g24637,g16586,g22884);
  AN2 AND2_3139(g19521,g513,g16739);
  AN2 AND2_3140(g22122,g6601,g19277);
  AN3 AND3_183(g12692,g10323,g3522,g3530);
  AN2 AND2_3141(g12761,g969,g7567);
  AN2 AND2_3142(g18284,g15071,g16164);
  AN2 AND2_3143(g16868,g5813,g14297);
  AN2 AND2_3144(g34497,g34275,g33072);
  AN2 AND2_3145(g28165,g27018,g22455);
  AN2 AND2_3146(g28523,g27704,g15585);
  AN2 AND2_3147(g18304,g1542,g16489);
  AN2 AND2_3148(g29182,g27163,g12730);
  AN2 AND2_3149(g29651,g2537,g29134);
  AN2 AND2_3150(g33412,g32362,g21411);
  AN4 AND4_194(I31322,g32921,g32922,g32923,g32924);
  AN2 AND2_3151(g16161,g5841,g14297);
  AN2 AND2_3152(g15611,g471,g13437);
  AN2 AND2_3153(g15722,g464,g13437);
  AN2 AND2_3154(g18622,g3480,g17062);
  AN2 AND2_3155(g22034,g5929,g19147);
  AN2 AND2_3156(g15080,g12855,g12983);
  AN2 AND2_3157(g18566,g2860,g16349);
  AN2 AND2_3158(g30126,g28582,g21058);
  AN2 AND2_3159(g14615,g10604,g10587);
  AN2 AND2_3160(g27214,g26026,g13901);
  AN2 AND2_3161(g34700,g34535,g20129);
  AN2 AND2_3162(g31229,g30288,g23949);
  AN3 AND3_184(g10720,g2704,g10219,g2689);
  AN2 AND2_3163(g21815,g3598,g20924);
  AN2 AND2_3164(g30250,g28744,g23939);
  AN2 AND2_3165(g27329,g12052,g26743);
  AN2 AND2_3166(g32309,g5160,g31528);
  AN2 AND2_3167(g27207,g26055,g16692);
  AN2 AND2_3168(g33896,g33314,g20771);
  AN2 AND2_3169(g31228,g20028,g29713);
  AN2 AND2_3170(g27539,g26576,g17745);
  AN2 AND2_3171(g29331,g29143,g22169);
  AN2 AND2_3172(g32224,g4300,g31327);
  AN2 AND2_3173(g34658,g34574,g18896);
  AN2 AND2_3174(g23187,g13989,g20010);
  AN2 AND2_3175(g26855,g2960,g24535);
  AN2 AND2_3176(g21975,g5523,g19074);
  AN2 AND2_3177(g27328,g12482,g26736);
  AN2 AND2_3178(g25089,g23317,g20553);
  AN2 AND2_3179(g32308,g31293,g23503);
  AN2 AND2_3180(g20215,g16479,g10476);
  AN2 AND2_3181(g29513,g28448,g14095);
  AN2 AND2_3182(g18139,g542,g17249);
  AN2 AND2_3183(g27538,g26549,g14744);
  AN2 AND2_3184(g18653,g4176,g16249);
  AN2 AND2_3185(g24501,g14000,g23182);
  AN2 AND2_3186(g24729,g22719,g23018);
  AN2 AND2_3187(g25088,g17601,g23491);
  AN2 AND2_3188(g17292,g1075,g13093);
  AN4 AND4_195(g11160,g6336,g7074,g6322,g10003);
  AN2 AND2_3189(g17153,g6311,g14943);
  AN3 AND3_185(I24033,g8219,g8443,g3747);
  AN2 AND2_3190(g18138,g546,g17249);
  AN4 AND4_196(I26531,g24099,g24100,g24101,g24102);
  AN2 AND2_3191(g21937,g5208,g18997);
  AN3 AND3_186(I17552,g13156,g11450,g11498);
  AN2 AND2_3192(g34338,g34099,g19905);
  AN2 AND2_3193(g24728,g16513,g23017);
  AN4 AND4_197(g16244,g11547,g11592,g6789,I17585);
  AN4 AND4_198(I31336,g31672,g31855,g32940,g32941);
  AN2 AND2_3194(g14035,g699,g11048);
  AN2 AND2_3195(g15650,g8362,g13413);
  AN2 AND2_3196(g34969,g34960,g19570);
  AN2 AND2_3197(g10684,g7998,g411);
  AN2 AND2_3198(g28703,g27925,g20680);
  AN2 AND2_3199(g18636,g3817,g17096);
  AN2 AND2_3200(g18415,g2108,g15373);
  AN2 AND2_3201(g31310,g30157,g27886);
  AN2 AND2_3202(g18333,g1691,g17873);
  AN2 AND2_3203(g30060,g29146,g10581);
  AN2 AND2_3204(g21791,g3368,g20391);
  AN2 AND2_3205(g28253,g23719,g27700);
  AN2 AND2_3206(g21884,g4104,g19801);
  AN2 AND2_3207(g11915,g1802,g7315);
  AN2 AND2_3208(g34968,g34952,g23203);
  AN2 AND2_3209(g23884,g4119,g19510);
  AN2 AND2_3210(g30197,g28661,g23859);
  AN2 AND2_3211(g31959,g4907,g30673);
  AN2 AND2_3212(g33379,g30984,g32364);
  AN4 AND4_199(g19462,g7850,g14182,g14177,g16646);
  AN2 AND2_3213(g25126,g16839,g23523);
  AN2 AND2_3214(g25987,g9501,g25015);
  AN4 AND4_200(I31017,g32480,g32481,g32482,g32483);
  AN2 AND2_3215(g13277,g3195,g11432);
  AN2 AND2_3216(g28236,g8515,g27971);
  AN2 AND2_3217(g34870,g34820,g19882);
  AN2 AND2_3218(g34527,g34303,g19603);
  AN2 AND2_3219(g24284,g4375,g22550);
  AN2 AND2_3220(g18664,g4332,g17367);
  AN2 AND2_3221(g27235,g25910,g19579);
  AN2 AND2_3222(g24304,g12875,g22228);
  AN2 AND2_3223(g26819,g106,g24490);
  AN2 AND2_3224(g27683,g25770,g23567);
  AN2 AND2_3225(g24622,g19856,g22866);
  AN3 AND3_187(g33742,g7828,g33142,I31600);
  AN2 AND2_3226(g26257,g4253,g25197);
  AN2 AND2_3227(g31944,g31745,g22146);
  AN2 AND2_3228(g11037,g6128,g9184);
  AN2 AND2_3229(g18576,g2868,g16349);
  AN2 AND2_3230(g18585,g2960,g16349);
  AN2 AND2_3231(g14193,g7178,g10590);
  AN2 AND2_3232(g18484,g2491,g15426);
  AN2 AND2_3233(g22109,g6455,g18833);
  AN2 AND2_3234(g32260,g31250,g20385);
  AN3 AND3_188(g28264,g7315,g1802,g27416);
  AN2 AND2_3235(g34503,g34278,g19437);
  AN2 AND2_3236(g34867,g34826,g20145);
  AN2 AND2_3237(g25969,g9310,g24987);
  AN2 AND2_3238(g18554,g2831,g15277);
  AN2 AND2_3239(g29620,g2399,g29097);
  AN2 AND2_3240(g33681,g33129,g7991);
  AN2 AND2_3241(g22108,g6439,g18833);
  AN2 AND2_3242(g18609,g3147,g16987);
  AN2 AND2_3243(g27414,g255,g26827);
  AN2 AND2_3244(g32195,g30734,g25451);
  AN2 AND2_3245(g24139,g17619,g21653);
  AN2 AND2_3246(g25968,g25215,g20739);
  AN2 AND2_3247(g18312,g1579,g16931);
  AN2 AND2_3248(g33802,g33097,g14545);
  AN2 AND2_3249(g33429,g32231,g29676);
  AN2 AND2_3250(g33857,g33267,g20445);
  AN2 AND2_3251(g29646,g1816,g28675);
  AN3 AND3_189(g30315,g29182,g7028,g5644);
  AN2 AND2_3252(g34581,g22864,g34312);
  AN2 AND2_3253(g18608,g15087,g16987);
  AN2 AND2_3254(g27407,g26488,g17522);
  AN2 AND2_3255(g18115,g460,g17015);
  AN4 AND4_201(I27534,g28039,g24128,g24129,g24130);
  AN4 AND4_202(g33730,g7202,g4621,g33127,g4633);
  AN2 AND2_3256(g32016,g8522,g31138);
  AN2 AND2_3257(g33428,g32230,g29672);
  AN2 AND2_3258(g34707,g34544,g20579);
  AN2 AND2_3259(g30202,g28667,g23863);
  AN2 AND2_3260(g25870,g24840,g16182);
  AN2 AND2_3261(g30257,g28750,g23952);
  AN3 AND3_190(g25411,g5062,g23764,I24546);
  AN2 AND2_3262(g26094,g24936,g9664);
  AN2 AND2_3263(g31765,g30128,g23968);
  AN2 AND2_3264(g24415,g4760,g22869);
  AN2 AND2_3265(g7763,g2965,g2960);
  AN2 AND2_3266(g24333,g4512,g22228);
  AN2 AND2_3267(g29369,g28209,g22341);
  AN2 AND2_3268(g14222,g8655,g11826);
  AN2 AND2_3269(g21922,g5112,g21468);
  AN2 AND2_3270(g22982,g19535,g19747);
  AN2 AND2_3271(g30111,g28565,g20917);
  AN2 AND2_3272(g18745,g5128,g17847);
  AN2 AND2_3273(g33690,g33146,g16280);
  AN2 AND2_3274(g30070,g29167,g9529);
  AN2 AND2_3275(g34111,g33733,g22936);
  AN2 AND2_3276(g18799,g6181,g15348);
  AN2 AND2_3277(g22091,g6415,g18833);
  AN2 AND2_3278(g23531,g10760,g18930);
  AN2 AND2_3279(g13853,g4549,g10620);
  AN2 AND2_3280(g18813,g6513,g15483);
  AN2 AND2_3281(g30590,g18911,g29812);
  AN2 AND2_3282(g21740,g3085,g20330);
  AN2 AND2_3283(g16599,g6601,g15030);
  AN2 AND2_3284(g26019,g5507,g25032);
  AN2 AND2_3285(g25503,g6888,g22529);
  AN2 AND2_3286(g18798,g6177,g15348);
  AN2 AND2_3287(g28542,g27405,g20275);
  AN2 AND2_3288(g31504,g29370,g10553);
  AN2 AND2_3289(g28453,g27582,g10233);
  AN2 AND2_3290(g27206,g26055,g16691);
  AN3 AND3_191(g33504,g32772,I31216,I31217);
  AN2 AND2_3291(g24664,g22652,g19741);
  AN2 AND2_3292(g29850,g28340,g24893);
  AN2 AND2_3293(g19911,g14707,g17748);
  AN2 AND2_3294(g34741,g8899,g34697);
  AN2 AND2_3295(g16598,g6283,g14899);
  AN2 AND2_3296(g15810,g3937,g14055);
  AN2 AND2_3297(g13524,g9995,g11910);
  AN2 AND2_3298(g17091,g8659,g12940);
  AN2 AND2_3299(g18184,g785,g17328);
  AN2 AND2_3300(g21953,g5377,g21514);
  AN2 AND2_3301(g18805,g6377,g15656);
  AN2 AND2_3302(g18674,g4340,g15758);
  AN2 AND2_3303(g23373,g13699,g20195);
  AN2 AND2_3304(g30094,g28544,g20767);
  AN4 AND4_203(g27759,g22457,g25224,g26424,g26213);
  AN2 AND2_3305(g25581,g19338,g24150);
  AN2 AND2_3306(g25450,g6888,g22497);
  AN2 AND2_3307(g32042,g27244,g31070);
  AN2 AND2_3308(g21800,g3546,g20924);
  AN2 AND2_3309(g24484,g16288,g23208);
  AN2 AND2_3310(g29896,g2599,g29171);
  AN2 AND2_3311(g27114,g25997,g16523);
  AN2 AND2_3312(g32255,g31248,g20381);
  AN2 AND2_3313(g31129,g1968,g30017);
  AN2 AND2_3314(g32189,g30824,g25369);
  AN2 AND2_3315(g21936,g5200,g18997);
  AN2 AND2_3316(g18732,g4961,g16877);
  AN2 AND2_3317(g27435,g26549,g17585);
  AN2 AND2_3318(g18934,g3133,g16096);
  AN2 AND2_3319(g30735,g29814,g22319);
  AN2 AND2_3320(g24554,g22490,g19541);
  AN2 AND2_3321(g27107,g26055,g16514);
  AN2 AND2_3322(g32270,g31254,g20444);
  AN2 AND2_3323(g16125,g5152,g14238);
  AN2 AND2_3324(g16532,g5252,g14841);
  AN2 AND2_3325(g25818,g8124,g24605);
  AN2 AND2_3326(g28530,g27383,g20240);
  AN2 AND2_3327(g31128,g12187,g30016);
  AN2 AND2_3328(g32188,g27586,g31376);
  AN2 AND2_3329(g25979,g24517,g19650);
  AN2 AND2_3330(g28346,g27243,g19800);
  AN2 AND2_3331(g7251,g452,g392);
  AN2 AND2_3332(g24312,g4501,g22228);
  AN2 AND2_3333(g18692,g4732,g16053);
  AN2 AND2_3334(g18761,g5471,g17929);
  AN2 AND2_3335(g33245,g32125,g19961);
  AN2 AND2_3336(g24608,g6500,g23425);
  AN2 AND2_3337(g25978,g9391,g25001);
  AN2 AND2_3338(g13313,g475,g11048);
  AN2 AND2_3339(g15967,g3913,g14058);
  AN2 AND2_3340(g30196,g28659,g23858);
  AN2 AND2_3341(g31323,g30150,g27907);
  AN2 AND2_3342(g29582,g27766,g28608);
  AN2 AND2_3343(g31299,g30123,g27800);
  AN2 AND2_3344(g17192,g1677,g13022);
  AN2 AND2_3345(g34196,g33682,g24485);
  AN2 AND2_3346(g21762,g3219,g20785);
  AN2 AND2_3347(g21964,g5441,g21514);
  AN2 AND2_3348(g25986,g5160,g25013);
  AN2 AND2_3349(g32030,g4172,g30937);
  AN2 AND2_3350(g24921,g23721,g20739);
  AN4 AND4_204(I31016,g30825,g31798,g32478,g32479);
  AN2 AND2_3351(g31298,g30169,g27886);
  AN2 AND2_3352(g34526,g34300,g19569);
  AN2 AND2_3353(g18400,g2012,g15373);
  AN2 AND2_3354(g10873,g3004,g9015);
  AN2 AND2_3355(g26077,g9607,g25233);
  AN2 AND2_3356(g24745,g650,g23550);
  AN2 AND2_3357(g29627,g28493,g11884);
  AN2 AND2_3358(g18214,g939,g15979);
  AN2 AND2_3359(g28292,g23781,g27762);
  AN2 AND2_3360(g29959,g28953,g12823);
  AN2 AND2_3361(g22862,g1570,g19673);
  AN3 AND3_192(g28153,g26424,g22763,g27031);
  AN2 AND2_3362(g18329,g1612,g17873);
  AN2 AND2_3363(g25067,g4722,g22885);
  AN2 AND2_3364(g25094,g23318,g20554);
  AN2 AND2_3365(g18207,g925,g15938);
  AN2 AND2_3366(g26689,g15754,g24431);
  AN2 AND2_3367(g29378,g28137,g22493);
  AN2 AND2_3368(g13808,g4543,g10607);
  AN2 AND2_3369(g18539,g2763,g15277);
  AN2 AND2_3370(g11036,g9806,g5774);
  AN2 AND2_3371(g26280,g13051,g25248);
  AN2 AND2_3372(g18328,g1657,g17873);
  AN2 AND2_3373(g27263,g25940,g19713);
  AN2 AND2_3374(g21909,g5041,g21468);
  AN2 AND2_3375(g31232,g30294,g23972);
  AN2 AND2_3376(g25150,g17480,g23547);
  AN2 AND2_3377(g22040,g5953,g19147);
  AN2 AND2_3378(g25801,g8097,g24585);
  AN2 AND2_3379(g26300,g1968,g25341);
  AN2 AND2_3380(g34866,g34819,g20106);
  AN2 AND2_3381(g28136,g27382,g23135);
  AN2 AND2_3382(g18538,g2759,g15277);
  AN2 AND2_3383(g15079,g2151,g12955);
  AN2 AND2_3384(g27332,g12538,g26758);
  AN2 AND2_3385(g29603,g2265,g29060);
  AN2 AND2_3386(g24674,g446,g23496);
  AN2 AND2_3387(g29742,g28288,g10233);
  AN2 AND2_3388(g21908,g5037,g21468);
  AN2 AND2_3389(g15078,g10361,g12955);
  AN2 AND2_3390(g33697,g33160,g13330);
  AN2 AND2_3391(g30001,g28490,g23486);
  AN2 AND2_3392(g31995,g28274,g30569);
  AN2 AND2_3393(g33856,g33266,g20442);
  AN2 AND2_3394(g26102,g1825,g25099);
  AN2 AND2_3395(g12135,g9684,g9959);
  AN2 AND2_3396(g31261,g14754,g30259);
  AN2 AND2_3397(g26157,g2093,g25136);
  AN2 AND2_3398(g27406,g26488,g17521);
  AN3 AND3_193(g34077,g22957,g9104,g33736);
  AN2 AND2_3399(g27962,g25954,g19597);
  AN2 AND2_3400(g27361,g26519,g17419);
  AN2 AND2_3401(g33880,g33290,g20568);
  AN4 AND4_205(I31042,g32515,g32516,g32517,g32518);
  AN2 AND2_3402(g18241,g1183,g16431);
  AN2 AND2_3403(g34706,g34496,g10570);
  AN2 AND2_3404(g21747,g3061,g20330);
  AN2 AND2_3405(g32160,g31001,g22995);
  AN2 AND2_3406(g30256,g28749,g23947);
  AN2 AND2_3407(g25526,g23720,g21400);
  AN2 AND2_3408(g28164,g8651,g27528);
  AN2 AND2_3409(g26231,g1854,g25300);
  AN3 AND3_194(g33512,g32830,I31256,I31257);
  AN2 AND2_3410(g14913,g1442,g10939);
  AN2 AND2_3411(g27500,g26400,g17672);
  AN2 AND2_3412(g29857,g28386,g23304);
  AN2 AND2_3413(g15817,g3921,g13929);
  AN2 AND2_3414(g14614,g11975,g11997);
  AN2 AND2_3415(g24761,g22751,g19852);
  AN2 AND2_3416(g19540,g1124,g15904);
  AN2 AND2_3417(g21814,g3594,g20924);
  AN2 AND2_3418(g18771,g5685,g15615);
  AN2 AND2_3419(g16023,g3813,g13584);
  AN2 AND2_3420(g16224,g14583,g14232);
  AN4 AND4_206(g11166,g8363,g269,g8296,I14225);
  AN2 AND2_3421(g18235,g1141,g16326);
  AN2 AND2_3422(g21751,g3167,g20785);
  AN2 AND2_3423(g21807,g3566,g20924);
  AN2 AND2_3424(g21772,g3259,g20785);
  AN2 AND2_3425(g26854,g2868,g24534);
  AN2 AND2_3426(g15783,g3215,g14098);
  AN2 AND2_3427(g21974,g5517,g19074);
  AN2 AND2_3428(g22062,g6093,g21611);
  AN2 AND2_3429(g18683,g4674,g15885);
  AN2 AND2_3430(g25866,g3853,g24648);
  AN2 AND2_3431(g24400,g3466,g23112);
  AN2 AND2_3432(g27221,g26055,g16747);
  AN3 AND3_195(g33831,g23088,g33149,g9104);
  AN2 AND2_3433(g28327,g27365,g19785);
  AN2 AND2_3434(g29549,g2012,g28900);
  AN2 AND2_3435(g34102,g33912,g23599);
  AN2 AND2_3436(g26511,g19265,g24364);
  AN2 AND2_3437(g34157,g33794,g20159);
  AN2 AND2_3438(g23639,g19050,g9104);
  AN4 AND4_207(I31267,g32840,g32841,g32842,g32843);
  AN2 AND2_3439(g10565,g8182,g424);
  AN2 AND2_3440(g28537,g6832,g27089);
  AN2 AND2_3441(g31499,g29801,g23446);
  AN3 AND3_196(g33499,g32737,I31191,I31192);
  AN2 AND2_3442(g14565,g11934,g11952);
  AN2 AND2_3443(g29548,g1798,g28575);
  AN2 AND2_3444(g23293,g9104,g19200);
  AN2 AND2_3445(g24329,g4462,g22228);
  AN2 AND2_3446(g30066,g28518,g20636);
  AN2 AND2_3447(g22851,g496,g19654);
  AN2 AND2_3448(g28108,g7975,g27237);
  AN2 AND2_3449(g30231,g28718,g23907);
  AN2 AND2_3450(g15823,g3945,g14116);
  AN2 AND2_3451(g34066,g33730,g19352);
  AN2 AND2_3452(g10034,g1521,g1500);
  AN2 AND2_3453(g25077,g23297,g20536);
  AN3 AND3_197(g33498,g32730,I31186,I31187);
  AN2 AND2_3454(g23265,g20069,g20132);
  AN2 AND2_3455(g24328,g4567,g22228);
  AN3 AND3_198(g28283,g7380,g2361,g27445);
  AN2 AND2_3456(g18515,g2643,g15509);
  AN2 AND2_3457(g23416,g20082,g20321);
  AN2 AND2_3458(g18414,g2102,g15373);
  AN2 AND2_3459(g31989,g31770,g22200);
  AN2 AND2_3460(g14641,g11994,g12020);
  AN3 AND3_199(g28303,g7462,g2629,g27494);
  AN2 AND2_3461(g27106,g26026,g16512);
  AN2 AND2_3462(g21841,g3857,g21070);
  AN2 AND2_3463(g21992,g5599,g19074);
  AN2 AND2_3464(g34876,g34844,g20534);
  AN2 AND2_3465(g18407,g2016,g15373);
  AN2 AND2_3466(g25923,g24443,g19443);
  AN2 AND2_3467(g31988,g31768,g22199);
  AN2 AND2_3468(g33722,g33175,g19445);
  AN2 AND2_3469(g33924,g33335,g33346);
  AN2 AND2_3470(g32419,g4955,g31000);
  AN2 AND2_3471(g15966,g3462,g13555);
  AN4 AND4_208(g28982,g27163,g12687,g20682,I27349);
  AN2 AND2_3472(g31271,g29706,g23300);
  AN2 AND2_3473(g12812,g518,g9158);
  AN2 AND2_3474(g34763,g34689,g19915);
  AN2 AND2_3475(g15631,g168,g13437);
  AN2 AND2_3476(g27033,g25767,g19273);
  AN2 AND2_3477(g27371,g26400,g17473);
  AN2 AND2_3478(g32418,g31126,g16239);
  AN2 AND2_3479(g26287,g2138,g25225);
  AN2 AND2_3480(g27234,g26055,g16814);
  AN2 AND2_3481(g25102,g4727,g22885);
  AN2 AND2_3482(g21835,g3802,g20453);
  AN2 AND2_3483(g32170,g31671,g27779);
  AN2 AND2_3484(g13567,g10102,g11948);
  AN2 AND2_3485(g22047,g6077,g21611);
  AN2 AND2_3486(g26307,g13070,g25288);
  AN2 AND2_3487(g26085,g11906,g25070);
  AN2 AND2_3488(g29626,g28584,g11415);
  AN3 AND3_200(g33461,g32463,I31001,I31002);
  AN2 AND2_3489(g16669,g5611,g14993);
  AN2 AND2_3490(g33342,g32226,g20660);
  AN3 AND3_201(g29323,g28539,g6905,g3639);
  AN2 AND2_3491(g23007,g681,g20248);
  AN2 AND2_3492(g31145,g9970,g30052);
  AN2 AND2_3493(g18441,g2246,g18008);
  AN2 AND2_3494(g18584,g2950,g16349);
  AN2 AND2_3495(g24771,g7028,g23605);
  AN2 AND2_3496(g18206,g918,g15938);
  AN2 AND2_3497(g29533,g28958,g22417);
  AN2 AND2_3498(g12795,g1312,g7601);
  AN2 AND2_3499(g16668,g5543,g14962);
  AN2 AND2_3500(g16842,g6279,g14861);
  AN2 AND2_3501(g17574,g9554,g14546);
  AN2 AND2_3502(g33887,g33298,g20615);
  AN2 AND2_3503(g18759,g5467,g17929);
  AN2 AND2_3504(g22051,g6105,g21611);
  AN2 AND2_3505(g22072,g6259,g19210);
  AN2 AND2_3506(g18725,g4912,g16077);
  AN2 AND2_3507(g32167,g3853,g31194);
  AN2 AND2_3508(g32194,g30601,g28436);
  AN2 AND2_3509(g25876,g3470,g24667);
  AN3 AND3_202(g33529,g32953,I31341,I31342);
  AN4 AND4_209(I31201,g31672,g31831,g32745,g32746);
  AN2 AND2_3510(g27507,g26549,g17683);
  AN4 AND4_210(I31277,g32856,g32857,g32858,g32859);
  AN2 AND2_3511(g18114,g452,g17015);
  AN2 AND2_3512(g28192,g8891,g27415);
  AN2 AND2_3513(g18758,g7004,g15595);
  AN2 AND2_3514(g31528,g19050,g29814);
  AN2 AND2_3515(g26341,g24746,g20105);
  AN2 AND2_3516(g18435,g2173,g18008);
  AN3 AND3_203(g33528,g32946,I31336,I31337);
  AN2 AND2_3517(g34287,g11370,g34124);
  AN2 AND2_3518(g19661,g5489,g16969);
  AN2 AND2_3519(g33843,g33256,g20325);
  AN2 AND2_3520(g21720,g376,g21037);
  AN2 AND2_3521(g33330,g32211,g20588);
  AN2 AND2_3522(g26156,g2028,g25135);
  AN2 AND2_3523(g18107,g429,g17015);
  AN4 AND4_211(g27421,g8038,g26314,g9187,g9077);
  AN3 AND3_204(g34085,g33761,g9104,g18957);
  AN2 AND2_3524(g28663,g27566,g20624);
  AN2 AND2_3525(g32401,g31116,g13432);
  AN2 AND2_3526(g34076,g33694,g19519);
  AN2 AND2_3527(g30596,g30279,g18947);
  AN2 AND2_3528(g26180,g2587,g25156);
  AN2 AND2_3529(g26670,g13385,g24428);
  AN2 AND2_3530(g21746,g3045,g20330);
  AN2 AND2_3531(g33365,g32267,g20994);
  AN2 AND2_3532(g32119,g31609,g29939);
  AN2 AND2_3533(g30243,g28731,g23929);
  AN2 AND2_3534(g31132,g29504,g22987);
  AN2 AND2_3535(g18744,g5124,g17847);
  AN2 AND2_3536(g34054,g33778,g22942);
  AN2 AND2_3537(g31960,g31749,g22153);
  AN2 AND2_3538(g33869,g33279,g20543);
  AN2 AND2_3539(g14537,g10550,g10529);
  AN2 AND2_3540(g18345,g1736,g17955);
  AN2 AND2_3541(g19715,g9679,g17120);
  AN4 AND4_212(I31037,g32508,g32509,g32510,g32511);
  AN2 AND2_3542(g29856,g28385,g23303);
  AN4 AND4_213(g17780,g6772,g11592,g11640,I18782);
  AN2 AND2_3543(g21465,g16155,g13663);
  AN2 AND2_3544(g18399,g2024,g15373);
  AN2 AND2_3545(g29880,g1936,g29149);
  AN2 AND2_3546(g33868,g33278,g20542);
  AN2 AND2_3547(g26839,g2988,g24516);
  AN2 AND2_3548(g27541,g26278,g23334);
  AN2 AND2_3549(g30269,g28778,g23970);
  AN2 AND2_3550(g22846,g9386,g20676);
  AN2 AND2_3551(g21983,g5555,g19074);
  AN2 AND2_3552(g28553,g27187,g10290);
  AN3 AND3_205(g25456,g5752,g22210,I24579);
  AN2 AND2_3553(g18398,g2020,g15373);
  AN2 AND2_3554(g29512,g2161,g28793);
  AN2 AND2_3555(g32313,g31303,g23515);
  AN4 AND4_214(I31352,g32963,g32964,g32965,g32966);
  AN2 AND2_3556(g21806,g3558,g20924);
  AN2 AND2_3557(g26838,g2860,g24515);
  AN2 AND2_3558(g18141,g568,g17533);
  AN2 AND2_3559(g30268,g28777,g23969);
  AN2 AND2_3560(g18652,g4172,g16249);
  AN2 AND2_3561(g18804,g15163,g15656);
  AN2 AND2_3562(g34341,g34101,g19952);
  AN2 AND2_3563(g25916,g24432,g19434);
  AN2 AND2_3564(g16610,g5260,g14918);
  AN2 AND2_3565(g16705,g6299,g15024);
  AN2 AND2_3566(g17152,g8635,g12997);
  AN2 AND2_3567(g31225,g30276,g21012);
  AN2 AND2_3568(g32276,g31646,g30313);
  AN4 AND4_215(g27724,g22417,g25208,g26424,g26190);
  AN2 AND2_3569(g34655,g34573,g18885);
  AN4 AND4_216(I31266,g31327,g31843,g32838,g32839);
  AN2 AND2_3570(g27359,g26488,g17416);
  AN2 AND2_3571(g30180,g28635,g23820);
  AN2 AND2_3572(g27325,g12478,g26724);
  AN2 AND2_3573(g30670,g11330,g29359);
  AN2 AND2_3574(g31471,g29754,g23399);
  AN2 AND2_3575(g32305,g31287,g20567);
  AN2 AND2_3576(g32053,g14176,g31509);
  AN3 AND3_206(g33471,g32535,I31051,I31052);
  AN2 AND2_3577(g34180,g33716,g24373);
  AN2 AND2_3578(g33087,g32391,g18888);
  AN2 AND2_3579(g18263,g1249,g16000);
  AN2 AND2_3580(g32254,g31247,g20379);
  AN2 AND2_3581(g27535,g26519,g17737);
  AN2 AND2_3582(g26487,g15702,g24359);
  AN2 AND2_3583(g27434,g26549,g17584);
  AN2 AND2_3584(g27358,g26400,g17415);
  AN2 AND2_3585(g25076,g12805,g23479);
  AN2 AND2_3586(g25085,g4912,g22908);
  AN2 AND2_3587(g18332,g1677,g17873);
  AN2 AND2_3588(g19784,g2775,g15877);
  AN2 AND2_3589(g28252,g27159,g19682);
  AN2 AND2_3590(g12920,g1227,g10960);
  AN2 AND2_3591(g18135,g136,g17249);
  AN2 AND2_3592(g34335,g8461,g34197);
  AN2 AND2_3593(g25054,g12778,g23452);
  AN2 AND2_3594(g24725,g19587,g23012);
  AN2 AND2_3595(g30930,g29915,g23342);
  AN2 AND2_3596(g32036,g31469,g13486);
  AN2 AND2_3597(g27121,g136,g26326);
  AN3 AND3_207(g29316,g28528,g6875,g3288);
  AN2 AND2_3598(g19354,g471,g16235);
  AN2 AND2_3599(g33244,g32190,g23152);
  AN2 AND2_3600(g32177,g30608,g25214);
  AN2 AND2_3601(g18406,g2060,g15373);
  AN2 AND2_3602(g13349,g4933,g11780);
  AN4 AND4_217(I31167,g32696,g32697,g32698,g32699);
  AN3 AND3_208(I18785,g13156,g6767,g11498);
  AN2 AND2_3603(g26279,g4249,g25213);
  AN2 AND2_3604(g18361,g1821,g17955);
  AN2 AND2_3605(g24758,g6523,g23733);
  AN2 AND2_3606(g23130,g728,g20248);
  AN2 AND2_3607(g34667,g34471,g33424);
  AN2 AND2_3608(g34694,g34530,g19885);
  AN2 AND2_3609(g17405,g1422,g13137);
  AN2 AND2_3610(g11083,g8836,g802);
  AN2 AND2_3611(g34965,g34949,g23084);
  AN2 AND2_3612(g30131,g28589,g21178);
  AN2 AND2_3613(g31069,g29793,g14150);
  AN2 AND2_3614(g19671,g1454,g16155);
  AN2 AND2_3615(g29989,g29006,g10489);
  AN2 AND2_3616(g18500,g2421,g15426);
  AN2 AND2_3617(g22020,g5863,g19147);
  AN2 AND2_3618(g27682,g25777,g23565);
  AN2 AND2_3619(g23165,g13954,g19964);
  AN2 AND2_3620(g28183,g27024,g19421);
  AN2 AND2_3621(g28673,g1373,g27122);
  AN2 AND2_3622(g33810,g33427,g12768);
  AN2 AND2_3623(g27291,g11969,g26653);
  AN2 AND2_3624(g29611,g28540,g14209);
  AN2 AND2_3625(g33657,g30991,g33443);
  AN2 AND2_3626(g26286,g2126,g25389);
  AN2 AND2_3627(g29988,g29187,g12235);
  AN2 AND2_3628(g29924,g13031,g29190);
  AN2 AND2_3629(g34487,g34416,g18983);
  AN2 AND2_3630(g13566,g7092,g12358);
  AN2 AND2_3631(g22046,g6073,g21611);
  AN2 AND2_3632(g26306,g13087,g25286);
  AN2 AND2_3633(g24849,g4165,g22227);
  AN2 AND2_3634(g33879,g33289,g20566);
  AN2 AND2_3635(g24940,g5011,g23971);
  AN2 AND2_3636(g24399,g3133,g23067);
  AN2 AND2_3637(g34502,g26363,g34343);
  AN2 AND2_3638(g30210,g28684,g23877);
  AN2 AND2_3639(g34557,g34352,g20555);
  AN2 AND2_3640(g23006,g19575,g19776);
  AN2 AND2_3641(g23475,g19070,g8971);
  AN2 AND2_3642(g33878,g33288,g20565);
  AN4 AND4_218(I31022,g32487,g32488,g32489,g32490);
  AN2 AND2_3643(g18221,g1018,g16100);
  AN2 AND2_3644(g22113,g6561,g19277);
  AN2 AND2_3645(g21863,g3957,g21070);
  AN2 AND2_3646(g26815,g4108,g24528);
  AN2 AND2_3647(g24141,g17657,g21656);
  AN2 AND2_3648(g34279,g34231,g19208);
  AN4 AND4_219(g11139,g5990,g7051,g5976,g9935);
  AN2 AND2_3649(g33886,g33297,g20614);
  AN2 AND2_3650(g27134,g25997,g16602);
  AN2 AND2_3651(g30278,g28818,g23988);
  AN2 AND2_3652(g27029,g26327,g11031);
  AN2 AND2_3653(g18613,g3338,g17200);
  AN2 AND2_3654(g31792,g30214,g24017);
  AN2 AND2_3655(g32166,g31007,g23029);
  AN2 AND2_3656(g32009,g31782,g22224);
  AN2 AND2_3657(g25993,g2610,g25025);
  AN2 AND2_3658(g31967,g31755,g22167);
  AN2 AND2_3659(g31994,g31775,g22215);
  AN2 AND2_3660(g22105,g6494,g18833);
  AN4 AND4_220(I31276,g31376,g31844,g32854,g32855);
  AN2 AND2_3661(g27028,g26342,g1157);
  AN2 AND2_3662(g29199,g27187,g12687);
  AN2 AND2_3663(g32008,g31781,g22223);
  AN2 AND2_3664(g25965,g2208,g24980);
  AN2 AND2_3665(g29650,g28949,g22472);
  AN2 AND2_3666(g29736,g28522,g10233);
  AN2 AND2_3667(g16160,g5499,g14262);
  AN2 AND2_3668(g29887,g28417,g23351);
  AN2 AND2_3669(g21703,g146,g20283);
  AN2 AND2_3670(g18273,g1287,g16031);
  AN2 AND2_3671(g24332,g4459,g22228);
  AN2 AND2_3672(g18106,g411,g17015);
  AN2 AND2_3673(g20135,g16258,g16695);
  AN2 AND2_3674(g18605,g3129,g16987);
  AN2 AND2_3675(g13415,g837,g11048);
  AN2 AND2_3676(g21347,g1339,g15750);
  AN2 AND2_3677(g13333,g4743,g11755);
  AN2 AND2_3678(g33425,g32380,g21466);
  AN2 AND2_3679(g28213,g27720,g23380);
  AN2 AND2_3680(g15679,g3470,g13555);
  AN2 AND2_3681(g18812,g6509,g15483);
  AN2 AND2_3682(g10948,g7880,g1478);
  AN2 AND2_3683(g18463,g2375,g15224);
  AN2 AND2_3684(g33919,g33438,g10795);
  AN2 AND2_3685(g24406,g13623,g22860);
  AN2 AND2_3686(g29528,g2429,g28874);
  AN4 AND4_221(I31036,g30673,g31802,g32506,g32507);
  AN2 AND2_3687(g24962,g23194,g20210);
  AN2 AND2_3688(g29843,g28373,g23289);
  AN2 AND2_3689(g21781,g3408,g20391);
  AN2 AND2_3690(g29330,g29114,g18894);
  AN2 AND2_3691(g16617,g6287,g14940);
  AN2 AND2_3692(g25502,g6946,g22527);
  AN2 AND2_3693(g15678,g1094,g13846);
  AN4 AND4_222(I31101,g30735,g31813,g32601,g32602);
  AN4 AND4_223(I31177,g32710,g32711,g32712,g32713);
  AN2 AND2_3694(g18951,g3484,g16124);
  AN2 AND2_3695(g30187,g28643,g23840);
  AN2 AND2_3696(g18371,g1870,g15171);
  AN3 AND3_209(g8721,g385,g376,g365);
  AN2 AND2_3697(g28205,g27516,g16746);
  AN2 AND2_3698(g18234,g1129,g16326);
  AN2 AND2_3699(g34187,g33708,g24397);
  AN2 AND2_3700(g17769,g1146,g13188);
  AN2 AND2_3701(g21952,g5366,g21514);
  AN2 AND2_3702(g28311,g9792,g27679);
  AN2 AND2_3703(g23372,g16448,g20194);
  AN2 AND2_3704(g29869,g2331,g29129);
  AN2 AND2_3705(g21821,g3723,g20453);
  AN2 AND2_3706(g17768,g13325,g10741);
  AN4 AND4_224(I26530,g26365,g24096,g24097,g24098);
  AN2 AND2_3707(g18795,g6163,g15348);
  AN2 AND2_3708(g30937,g22626,g29814);
  AN2 AND2_3709(g29868,g2227,g29128);
  AN2 AND2_3710(g27649,g10820,g25820);
  AN2 AND2_3711(g34143,g33934,g23828);
  AN2 AND2_3712(g16595,g5921,g14697);
  AN2 AND2_3713(g21790,g3454,g20391);
  AN2 AND2_3714(g24004,g37,g21225);
  AN2 AND2_3715(g33086,g32390,g18887);
  AN2 AND2_3716(g27648,g25882,g8974);
  AN2 AND2_3717(g24221,g232,g22594);
  AN2 AND2_3718(g27491,g26576,g17652);
  AN2 AND2_3719(g26486,g4423,g24358);
  AN2 AND2_3720(g18514,g2629,g15509);
  AN2 AND2_3721(g29709,g2116,g29121);
  AN2 AND2_3722(g34169,g33804,g31227);
  AN2 AND2_3723(g21873,g6946,g19801);
  AN2 AND2_3724(g18507,g2595,g15509);
  AN2 AND2_3725(g22027,g5889,g19147);
  AN2 AND2_3726(g23873,g21222,g10815);
  AN2 AND2_3727(g15875,g3961,g13963);
  AN2 AND2_3728(g30168,g28623,g23794);
  AN2 AND2_3729(g29708,g1955,g29082);
  AN2 AND2_3730(g33817,g33235,g20102);
  AN2 AND2_3731(g11115,g6133,g9954);
  AN2 AND2_3732(g33322,g32202,g20450);
  AN2 AND2_3733(g34410,g34204,g21427);
  AN2 AND2_3734(g27981,g26751,g23924);
  AN2 AND2_3735(g25815,g8155,g24603);
  AN2 AND2_3736(g31125,g29502,g22973);
  AN2 AND2_3737(g32176,g2779,g31623);
  AN4 AND4_225(I31166,g30673,g31825,g32694,g32695);
  AN4 AND4_226(g26223,g24688,g10678,g10658,g8757);
  AN2 AND2_3738(g31977,g31764,g22179);
  AN3 AND3_210(g33532,g32974,I31356,I31357);
  AN2 AND2_3739(g33901,g33317,g20920);
  AN2 AND2_3740(g34479,g34403,g18905);
  AN2 AND2_3741(g34666,g34587,g19144);
  AN2 AND2_3742(g25187,g12296,g23629);
  AN2 AND2_3743(g18163,g79,g17433);
  AN2 AND2_3744(g15837,g3255,g14127);
  AN2 AND2_3745(g32154,g31277,g14184);
  AN2 AND2_3746(g34363,g34148,g20389);
  AN2 AND2_3747(g25975,g9434,g24999);
  AN2 AND2_3748(g34217,g33736,g22876);
  AN2 AND2_3749(g22710,g19358,g19600);
  AN2 AND2_3750(g30015,g29040,g10519);
  AN2 AND2_3751(g21834,g3752,g20453);
  AN2 AND2_3752(g22003,g5736,g21562);
  AN2 AND2_3753(g34478,g34402,g18904);
  AN2 AND2_3754(g28152,g26297,g27279);
  AN2 AND2_3755(g26084,g24926,g9602);
  AN4 AND4_227(g28846,g21434,g26424,g25399,g27474);
  AN2 AND2_3756(g24812,g19662,g22192);
  AN2 AND2_3757(g19855,g2787,g15962);
  AN2 AND2_3758(g33353,g32240,g20732);
  AN2 AND2_3759(g25143,g4922,g22908);
  AN2 AND2_3760(g34486,g34412,g18953);
  AN2 AND2_3761(g18541,g2767,g15277);
  AN4 AND4_228(g27395,g8046,g26314,g9187,g9077);
  AN2 AND2_3762(g33680,g33128,g4688);
  AN2 AND2_3763(g18473,g2342,g15224);
  AN2 AND2_3764(g27262,g25997,g17092);
  AN2 AND2_3765(g26179,g2504,g25155);
  AN2 AND2_3766(g12794,g1008,g7567);
  AN3 AND3_211(I17529,g13156,g11450,g6756);
  AN2 AND2_3767(g34556,g34350,g20537);
  AN2 AND2_3768(g18789,g6035,g15634);
  AN2 AND2_3769(g21453,g16713,g13625);
  AN2 AND2_3770(g22081,g6279,g19210);
  AN2 AND2_3771(g29602,g2020,g28962);
  AN2 AND2_3772(g29810,g28259,g11317);
  AN2 AND2_3773(g29774,g28287,g10233);
  AN2 AND2_3774(g34580,g29539,g34311);
  AN2 AND2_3775(g26178,g2389,g25473);
  AN4 AND4_229(g16194,g11547,g6782,g11640,I17529);
  AN2 AND2_3776(g27633,g13076,g25766);
  AN2 AND2_3777(g21913,g5069,g21468);
  AN2 AND2_3778(g29375,g13946,g28370);
  AN2 AND2_3779(g30223,g28702,g23895);
  AN4 AND4_230(g13805,g11489,g11394,g11356,I16129);
  AN2 AND2_3780(g18788,g6031,g15634);
  AN2 AND2_3781(g18724,g4907,g16077);
  AN2 AND2_3782(g25884,g11153,g24711);
  AN2 AND2_3783(g18359,g1825,g17955);
  AN2 AND2_3784(g34223,g33744,g22876);
  AN2 AND2_3785(g18325,g1624,g17873);
  AN2 AND2_3786(g26186,g24580,g23031);
  AN2 AND2_3787(g23436,g676,g20375);
  AN2 AND2_3788(g18535,g2741,g15277);
  AN2 AND2_3789(g18434,g2217,g18008);
  AN2 AND2_3790(g18358,g1811,g17955);
  AN2 AND2_3791(g31966,g31754,g22166);
  AN2 AND2_3792(g30084,g28534,g20700);
  AN2 AND2_3793(g27521,g26519,g14700);
  AN2 AND2_3794(g29337,g29166,g22180);
  AN2 AND2_3795(g17786,g1489,g13216);
  AN2 AND2_3796(g30110,g28564,g20916);
  AN2 AND2_3797(g25479,g22646,g9917);
  AN2 AND2_3798(g34084,g9214,g33851);
  AN2 AND2_3799(g15075,g12850,g12955);
  AN2 AND2_3800(g31017,g29479,g22841);
  AN2 AND2_3801(g34110,g33732,g22935);
  AN2 AND2_3802(g25217,g12418,g23698);
  AN2 AND2_3803(g33364,g32264,g20921);
  AN2 AND2_3804(g18121,g424,g17015);
  AN2 AND2_3805(g22090,g6404,g18833);
  AN2 AND2_3806(g30179,g28634,g23819);
  AN2 AND2_3807(g24507,g22304,g19429);
  AN2 AND2_3808(g18344,g1740,g17955);
  AN3 AND3_212(g19581,g15843,g1500,g10918);
  AN2 AND2_3809(g34179,g33686,g24372);
  AN4 AND4_231(g27440,g8046,g26314,g518,g504);
  AN2 AND2_3810(g21464,g16181,g10872);
  AN4 AND4_232(g28020,g23032,g26241,g26424,g25542);
  AN2 AND2_3811(g28583,g12009,g27112);
  AN2 AND2_3812(g30178,g28632,g23815);
  AN2 AND2_3813(g9479,g305,g324);
  AN2 AND2_3814(g24421,g3835,g23139);
  AN2 AND2_3815(g34178,g33712,g24361);
  AN2 AND2_3816(g34740,g34664,g19414);
  AN2 AND2_3817(g16616,g6267,g14741);
  AN4 AND4_233(g10756,g3990,g6928,g3976,g8595);
  AN2 AND2_3818(g18682,g4646,g15885);
  AN4 AND4_234(I31176,g31579,g31827,g32708,g32709);
  AN2 AND2_3819(g30186,g28641,g23839);
  AN2 AND2_3820(g27247,g2759,g26745);
  AN4 AND4_235(I31092,g32589,g32590,g32591,g32592);
  AN2 AND2_3821(g18291,g1437,g16449);
  AN2 AND2_3822(g24012,g14496,g21561);
  AN2 AND2_3823(g17182,g8579,g13016);
  AN2 AND2_3824(g21797,g3518,g20924);
  AN2 AND2_3825(g34186,g33705,g24396);
  AN2 AND2_3826(g34685,g14164,g34550);
  AN2 AND2_3827(g25580,g19268,g24149);
  AN2 AND2_3828(g18173,g736,g17328);
  AN2 AND2_3829(g27389,g26519,g17503);
  AN2 AND2_3830(g34953,g34935,g19957);
  AN4 AND4_236(g27045,g10295,g3171,g3179,g26244);
  AN2 AND2_3831(g31309,g30132,g27837);
  AN4 AND4_237(I24699,g21127,g24054,g24055,g24056);
  AN2 AND2_3832(g32083,g947,g30735);
  AN2 AND2_3833(g32348,g2145,g31672);
  AN2 AND2_3834(g23292,g19879,g16726);
  AN2 AND2_3835(g25223,g22523,g10652);
  AN2 AND2_3836(g16704,g5957,g15018);
  AN2 AND2_3837(g27612,g25887,g8844);
  AN2 AND2_3838(g31224,g30280,g23932);
  AN2 AND2_3839(g32284,g31260,g20507);
  AN2 AND2_3840(g28113,g8016,g27242);
  AN2 AND2_3841(g26423,g19488,g24356);
  AN2 AND2_3842(g27099,g14094,g26352);
  AN2 AND2_3843(g15822,g3925,g13960);
  AN2 AND2_3844(g27388,g26519,g17502);
  AN2 AND2_3845(g27324,g10150,g26720);
  AN2 AND2_3846(g24541,g22626,g10851);
  AN2 AND2_3847(g32304,g31284,g20564);
  AN2 AND2_3848(g30936,g8830,g29916);
  AN2 AND2_3849(g28282,g23762,g27727);
  AN2 AND2_3850(g12099,g9619,g9888);
  AN2 AND2_3851(g27534,g26488,g17735);
  AN2 AND2_3852(g27098,g25868,g22528);
  AN2 AND2_3853(g28302,g23809,g27817);
  AN2 AND2_3854(g25084,g4737,g22885);
  AN2 AND2_3855(g27251,g26721,g26694);
  AN2 AND2_3856(g27272,g26055,g17144);
  AN2 AND2_3857(g25110,g10427,g23509);
  AN2 AND2_3858(g16808,g6653,g14825);
  AN2 AND2_3859(g19384,g667,g16310);
  AN2 AND2_3860(g18760,g5462,g17929);
  AN2 AND2_3861(g18134,g534,g17249);
  AN2 AND2_3862(g25922,g24959,g20065);
  AN2 AND2_3863(g34334,g34090,g19865);
  AN2 AND2_3864(g24788,g11384,g23111);
  AN2 AND2_3865(g31495,g1913,g30309);
  AN2 AND2_3866(g24724,g17624,g22432);
  AN2 AND2_3867(g29599,g1710,g29018);
  AN3 AND3_213(g33495,g32707,I31171,I31172);
  AN2 AND2_3868(g22717,g9291,g20212);
  AN2 AND2_3869(g16177,g5128,g14238);
  AN2 AND2_3870(g24325,g4543,g22228);
  AN2 AND2_3871(g25179,g16928,g23611);
  AN2 AND2_3872(g26543,g12910,g24377);
  AN4 AND4_238(I27503,g19890,g24075,g24076,g28032);
  AN2 AND2_3873(g18506,g2571,g15509);
  AN2 AND2_3874(g22026,g5913,g19147);
  AN2 AND2_3875(g27462,g26576,g17612);
  AN2 AND2_3876(g33816,g33234,g20096);
  AN2 AND2_3877(g29598,g28823,g22342);
  AN2 AND2_3878(g16642,g6633,g14981);
  AN2 AND2_3879(g25178,g20241,g23608);
  AN2 AND2_3880(g15589,g411,g13334);
  AN2 AND2_3881(g32139,g31601,g29960);
  AN4 AND4_239(g27032,g7704,g5180,g5188,g26200);
  AN2 AND2_3882(g34964,g34947,g23060);
  AN2 AND2_3883(g33687,g33132,g4878);
  AN2 AND2_3884(g31976,g31762,g22178);
  AN2 AND2_3885(g31985,g4722,g30614);
  AN2 AND2_3886(g19735,g9740,g17135);
  AN2 AND2_3887(g27140,g25885,g22593);
  AN2 AND2_3888(g30216,g28691,g23882);
  AN2 AND2_3889(g27997,g26813,g23995);
  AN4 AND4_240(g28768,g21434,g26424,g25308,g27421);
  AN2 AND2_3890(g15836,g3187,g14104);
  AN2 AND2_3891(g31752,g30104,g23928);
  AN2 AND2_3892(g34216,g33778,g22689);
  AN2 AND2_3893(g31374,g29748,g23390);
  AN3 AND3_214(g29322,g29192,g7074,g6336);
  AN2 AND2_3894(g33374,g32289,g21221);
  AN2 AND2_3895(g16733,g5893,g14889);
  AN3 AND3_215(I18671,g13156,g11450,g6756);
  AN2 AND2_3896(g29532,g1878,g28861);
  AN2 AND2_3897(g29901,g28429,g23376);
  AN2 AND2_3898(g32333,g31326,g23559);
  AN2 AND2_3899(g15119,g4249,g14454);
  AN2 AND2_3900(g20682,g16238,g4646);
  AN4 AND4_241(g13771,g11441,g11355,g11302,I16111);
  AN3 AND3_216(g25417,g5712,g23816,I24552);
  AN2 AND2_3901(g23474,g13830,g20533);
  AN2 AND2_3902(g24682,g22662,g19754);
  AN2 AND2_3903(g22149,g14581,g18880);
  AN2 AND2_3904(g29783,g28329,g23246);
  AN2 AND2_3905(g21711,g291,g20283);
  AN2 AND2_3906(g26123,g1696,g25382);
  AN2 AND2_3907(g15118,g4253,g14454);
  AN2 AND2_3908(g34909,g34856,g20130);
  AN2 AND2_3909(g24291,g18660,g22550);
  AN2 AND2_3910(g30000,g23685,g29029);
  AN2 AND2_3911(g29656,g28515,g11666);
  AN2 AND2_3912(g34117,g33742,g19755);
  AN2 AND2_3913(g15749,g1454,g13273);
  AN2 AND2_3914(g18649,g4049,g17271);
  AN2 AND2_3915(g22097,g6451,g18833);
  AN2 AND2_3916(g27360,g26488,g17417);
  AN2 AND2_3917(g33842,g33255,g20322);
  AN2 AND2_3918(g18240,g15066,g16431);
  AN2 AND2_3919(g22104,g6444,g18833);
  AN2 AND2_3920(g17149,g232,g13255);
  AN2 AND2_3921(g33392,g32344,g21362);
  AN2 AND2_3922(g18648,g4045,g17271);
  AN2 AND2_3923(g18491,g2518,g15426);
  AN2 AND2_3924(g31489,g2204,g30305);
  AN2 AND2_3925(g26230,g1768,g25385);
  AN2 AND2_3926(g25964,g1783,g24979);
  AN3 AND3_217(g33489,g32665,I31141,I31142);
  AN2 AND2_3927(g21606,g15959,g13763);
  AN3 AND3_218(g27162,g26171,g8259,g2208);
  AN2 AND2_3928(g34568,g34379,g17512);
  AN2 AND2_3929(g34747,g34671,g19527);
  AN2 AND2_3930(g23606,g16927,g20679);
  AN2 AND2_3931(g29336,g4704,g28363);
  AN2 AND2_3932(g15704,g3440,g13504);
  AN2 AND2_3933(g30242,g28730,g23927);
  AN2 AND2_3934(g18604,g3125,g16987);
  AN2 AND2_3935(g21303,g10120,g17625);
  AN2 AND2_3936(g16485,g5563,g14924);
  AN2 AND2_3937(g18755,g5343,g15595);
  AN2 AND2_3938(g31525,g29892,g23526);
  AN2 AND2_3939(g31488,g1779,g30302);
  AN2 AND2_3940(g31016,g29478,g22840);
  AN3 AND3_219(g33525,g32925,I31321,I31322);
  AN3 AND3_220(g33488,g32658,I31136,I31137);
  AN2 AND2_3941(g28249,g27152,g19677);
  AN2 AND2_3942(g15809,g3917,g14154);
  AN2 AND2_3943(g18770,g15153,g15615);
  AN3 AND3_221(g22369,g9354,g7717,g20783);
  AN2 AND2_3944(g18563,g2890,g16349);
  AN2 AND2_3945(g18981,g11206,g16158);
  AN2 AND2_3946(g21750,g3161,g20785);
  AN2 AND2_3947(g28248,g27150,g19676);
  AN2 AND2_3948(g29966,g23617,g28970);
  AN2 AND2_3949(g28710,g27589,g20703);
  AN2 AND2_3950(g15808,g3590,g14048);
  AN2 AND2_3951(g21982,g5547,g19074);
  AN2 AND2_3952(g27451,g26400,g17599);
  AN2 AND2_3953(g26391,g19593,g25555);
  AN3 AND3_222(I26948,g24981,g26424,g22698);
  AN2 AND2_3954(g23381,g7239,g21413);
  AN2 AND2_3955(g27220,g26026,g16743);
  AN2 AND2_3956(g33830,g33382,g20166);
  AN2 AND2_3957(g29631,g1682,g28656);
  AN2 AND2_3958(g32312,g31302,g20591);
  AN2 AND2_3959(g32200,g27468,g31376);
  AN2 AND2_3960(g33893,g33313,g20706);
  AN2 AND2_3961(g28204,g26098,g27654);
  AN2 AND2_3962(g27628,g26400,g18061);
  AN2 AND2_3963(g34751,g34674,g19543);
  AN2 AND2_3964(g29364,g27400,g28321);
  AN2 AND2_3965(g10827,g8914,g4258);
  AN2 AND2_3966(g25909,g8745,g24875);
  AN2 AND2_3967(g32115,g31631,g29928);
  AN2 AND2_3968(g25543,g23795,g21461);
  AN2 AND2_3969(g12220,g1521,g7535);
  AN2 AND2_3970(g27246,g26690,g26673);
  AN2 AND2_3971(g33865,g33275,g20526);
  AN2 AND2_3972(g21796,g3512,g20924);
  AN2 AND2_3973(g30230,g28717,g23906);
  AN2 AND2_3974(g25908,g24782,g22520);
  AN2 AND2_3975(g18767,g15150,g17929);
  AN2 AND2_3976(g18794,g6154,g15348);
  AN2 AND2_3977(g34230,g33761,g22942);
  AN2 AND2_3978(g18395,g12849,g15373);
  AN2 AND2_3979(g32052,g31507,g13885);
  AN2 AND2_3980(g18262,g1259,g16000);
  AN2 AND2_3981(g22133,g6649,g19277);
  AN2 AND2_3982(g25569,I24684,I24685);
  AN2 AND2_3983(g21840,g15099,g21070);
  AN2 AND2_3984(g25568,I24679,I24680);
  AN2 AND2_3985(g18633,g6905,g17226);
  AN2 AND2_3986(g17133,g10683,g13222);
  AN2 AND2_3987(g34841,g34761,g20080);
  AN2 AND2_3988(g18191,g827,g17821);
  AN2 AND2_3989(g18719,g4894,g16795);
  AN2 AND2_3990(g22011,g15154,g21562);
  AN2 AND2_3991(g15874,g3893,g14079);
  AN2 AND2_3992(g24649,g6527,g23733);
  AN2 AND2_3993(g29571,g28452,g11762);
  AN2 AND2_3994(g11114,g5689,g10160);
  AN2 AND2_3995(g31270,g29692,g23282);
  AN2 AND2_3996(g16519,g5591,g14804);
  AN2 AND2_3997(g16176,g14596,g11779);
  AN2 AND2_3998(g16185,g3263,g14011);
  AN2 AND2_3999(g25123,g4732,g22885);
  AN2 AND2_4000(g18718,g4854,g15915);
  AN2 AND2_4001(g15693,g269,g13474);
  AN2 AND2_4002(g18521,g2667,g15509);
  AN2 AND2_4003(g31188,g20028,g29653);
  AN2 AND2_4004(g25814,g24760,g13323);
  AN2 AND2_4005(g27370,g26400,g17472);
  AN2 AND2_4006(g31124,g2259,g29997);
  AN2 AND2_4007(g32184,g30611,g25249);
  AN4 AND4_242(g28998,g17424,g25212,g26424,g27474);
  AN2 AND2_4008(g33124,g8945,g32296);
  AN3 AND3_223(g33678,g33149,g10710,g22319);
  AN2 AND2_4009(g24491,g10727,g22332);
  AN2 AND2_4010(g24903,g128,g23889);
  AN2 AND2_4011(g28233,g27827,g23411);
  AN2 AND2_4012(g16518,g5571,g14956);
  AN2 AND2_4013(g28182,g8770,g27349);
  AN2 AND2_4014(g25772,g24944,g24934);
  AN2 AND2_4015(g28672,g7577,g27017);
  AN2 AND2_4016(g24755,g16022,g23030);
  AN2 AND2_4017(g27151,g26026,g16626);
  AN2 AND2_4018(g34578,g24578,g34308);
  AN2 AND2_4019(g16637,g5949,g14968);
  AN2 AND2_4020(g22310,g19662,g20235);
  AN2 AND2_4021(g18440,g2255,g18008);
  AN2 AND2_4022(g13345,g4754,g11773);
  AN2 AND2_4023(g26275,g2417,g25349);
  AN2 AND2_4024(g30007,g29141,g12929);
  AN3 AND3_224(I24546,g5046,g5052,g9716);
  AN2 AND2_4025(g34586,g11025,g34317);
  AN2 AND2_4026(g18573,g2898,g16349);
  AN2 AND2_4027(g29687,g2407,g29097);
  AN2 AND2_4028(g22112,g6555,g19277);
  AN2 AND2_4029(g18247,g1178,g16431);
  AN2 AND2_4030(g29985,g28127,g20532);
  AN2 AND2_4031(g10890,g7858,g1105);
  AN2 AND2_4032(g21862,g3953,g21070);
  AN2 AND2_4033(g22050,g6088,g21611);
  AN2 AND2_4034(g23553,g19413,g11875);
  AN2 AND2_4035(g18389,g1974,g15171);
  AN2 AND2_4036(g29752,g28516,g10233);
  AN4 AND4_243(I31312,g32905,g32906,g32907,g32908);
  AN2 AND2_4037(g29954,g2299,g28796);
  AN2 AND2_4038(g21949,g5264,g18997);
  AN2 AND2_4039(g15712,g3791,g13521);
  AN2 AND2_4040(g18612,g3329,g17200);
  AN2 AND2_4041(g15914,g3905,g14024);
  AN2 AND2_4042(g25992,g2485,g25024);
  AN2 AND2_4043(g18388,g1968,g15171);
  AN2 AND2_4044(g19660,g12001,g16968);
  AN2 AND2_4045(g18324,g1644,g17873);
  AN2 AND2_4046(g24794,g11414,g23138);
  AN2 AND2_4047(g31219,g30265,g20875);
  AN2 AND2_4048(g34116,g33933,g25140);
  AN2 AND2_4049(g24395,g4704,g22845);
  AN3 AND3_225(g25510,g6444,g22300,I24619);
  AN2 AND2_4050(g18701,g4771,g16856);
  AN2 AND2_4051(g26684,g25407,g20673);
  AN2 AND2_4052(g21948,g5260,g18997);
  AN2 AND2_4053(g22096,g6434,g18833);
  AN2 AND2_4054(g32400,g4743,g30989);
  AN2 AND2_4055(g18777,g5808,g18065);
  AN2 AND2_4056(g18534,g2735,g15277);
  AN4 AND4_244(I14198,g225,g8237,g232,g8180);
  AN2 AND2_4057(g32013,g8673,g30614);
  AN2 AND2_4058(g30041,g28511,g23518);
  AN4 AND4_245(I31052,g32531,g32532,g32533,g32534);
  AN2 AND2_4059(g18251,g996,g16897);
  AN2 AND2_4060(g21702,g157,g20283);
  AN2 AND2_4061(g31218,g30271,g23909);
  AN2 AND2_4062(g16729,g5240,g14720);
  AN2 AND2_4063(g18272,g1283,g16031);
  AN2 AND2_4064(g21757,g3187,g20785);
  AN2 AND2_4065(g25579,g19422,g24147);
  AN2 AND2_4066(g30275,g28816,g23984);
  AN4 AND4_246(I24700,g24057,g24058,g24059,g24060);
  AN2 AND2_4067(g27227,g26026,g16771);
  AN2 AND2_4068(g33837,g33251,g20233);
  AN3 AND3_226(I24625,g6428,g6434,g10014);
  AN2 AND2_4069(g32207,g31221,g23323);
  AN2 AND2_4070(g26517,g15708,g24367);
  AN2 AND2_4071(g34746,g34670,g19526);
  AN2 AND2_4072(g34493,g34273,g19360);
  AN2 AND2_4073(g25578,g19402,g24146);
  AN2 AND2_4074(g15567,g392,g13312);
  AN2 AND2_4075(g27025,g26334,g7917);
  AN2 AND2_4076(g24191,g319,g22722);
  AN2 AND2_4077(g24719,g681,g23530);
  AN2 AND2_4078(g18462,g2361,g15224);
  AN2 AND2_4079(g25014,g17474,g23420);
  AN2 AND2_4080(g32328,g5853,g31554);
  AN2 AND2_4081(g29668,g28527,g14255);
  AN2 AND2_4082(g29842,g28372,g23284);
  AN2 AND2_4083(g27540,g26576,g17746);
  AN2 AND2_4084(g23564,g16882,g20648);
  AN4 AND4_247(g27058,g10323,g3522,g3530,g26264);
  AN2 AND2_4085(g30035,g22539,g28120);
  AN2 AND2_4086(g18140,g559,g17533);
  AN2 AND2_4087(g34340,g34100,g19950);
  AN2 AND2_4088(g27203,g26026,g16688);
  AN2 AND2_4089(g19596,g1094,g16681);
  AN2 AND2_4090(g26130,g24890,g19772);
  AN2 AND2_4091(g29525,g2169,g28837);
  AN2 AND2_4092(g21847,g3905,g21070);
  AN2 AND2_4093(g34684,g14178,g34545);
  AN2 AND2_4094(g10999,g7880,g1472);
  AN2 AND2_4095(g13833,g4546,g10613);
  AN3 AND3_227(I18819,g13156,g11450,g11498);
  AN2 AND2_4096(g26362,g19557,g25538);
  AN4 AND4_248(g27044,g7766,g5873,g5881,g26241);
  AN2 AND2_4097(g31470,g29753,g23398);
  AN2 AND2_4098(g23397,g11154,g20239);
  AN3 AND3_228(g33470,g32528,I31046,I31047);
  AN2 AND2_4099(g33915,g33140,g7846);
  AN2 AND2_4100(g32241,g31244,g20323);
  AN2 AND2_4101(g26165,g11980,g25153);
  AN4 AND4_249(g17793,g6772,g11592,g6789,I18803);
  AN4 AND4_250(g10998,g8567,g8509,g8451,g7650);
  AN2 AND2_4102(g18766,g5495,g17929);
  AN2 AND2_4103(g13048,g8558,g11043);
  AN2 AND2_4104(g23062,g718,g20248);
  AN2 AND2_4105(g27281,g9830,g26615);
  AN3 AND3_229(g24861,g3712,g23582,I24033);
  AN2 AND2_4106(g24573,g17198,g23716);
  AN2 AND2_4107(g34517,g34290,g19493);
  AN2 AND2_4108(g28148,g27355,g26093);
  AN2 AND2_4109(g14233,g8639,g11855);
  AN2 AND2_4110(g21933,g5212,g18997);
  AN2 AND2_4111(g27301,g11992,g26679);
  AN4 AND4_251(I14225,g8457,g255,g8406,g262);
  AN2 AND2_4112(g27957,g25947,g15995);
  AN2 AND2_4113(g7804,g2975,g2970);
  AN2 AND2_4114(g25041,g23261,g20494);
  AN2 AND2_4115(g13221,g6946,g11425);
  AN2 AND2_4116(g27120,g25878,g22543);
  AN4 AND4_252(g17690,g11547,g11592,g11640,I18671);
  AN2 AND2_4117(g29865,g1802,g29115);
  AN2 AND2_4118(g21851,g3901,g21070);
  AN2 AND2_4119(g21872,g4098,g19801);
  AN2 AND2_4120(g23872,g19389,g4157);
  AN2 AND2_4121(g15883,g9180,g14258);
  AN2 AND2_4122(g18360,g1830,g17955);
  AN2 AND2_4123(g31467,g30162,g27937);
  AN2 AND2_4124(g31494,g29792,g23435);
  AN2 AND2_4125(g28343,g27380,g19799);
  AN3 AND3_230(I24527,g9672,g9264,g5401);
  AN2 AND2_4126(g19655,g2729,g16966);
  AN3 AND3_231(g33467,g32505,I31031,I31032);
  AN3 AND3_232(g33494,g32700,I31166,I31167);
  AN2 AND2_4127(g24324,g4540,g22228);
  AN3 AND3_233(g27146,g26148,g8187,g1648);
  AN2 AND2_4128(g27645,g26488,g15344);
  AN2 AND2_4129(g26863,g24974,g24957);
  AN2 AND2_4130(g18447,g2208,g18008);
  AN2 AND2_4131(g30193,g28650,g23848);
  AN2 AND2_4132(g24777,g11345,g23066);
  AN2 AND2_4133(g27699,g26396,g20766);
  AN2 AND2_4134(g16653,g8343,g13850);
  AN2 AND2_4135(g18162,g686,g17433);
  AN2 AND2_4136(g25983,g2476,g25009);
  AN2 AND2_4137(g29610,g28483,g8026);
  AN2 AND2_4138(g30165,g28619,g23788);
  AN2 AND2_4139(g22129,g6633,g19277);
  AN2 AND2_4140(g34523,g9162,g34351);
  AN2 AND2_4141(g22002,g5706,g21562);
  AN2 AND2_4142(g22057,g15159,g21611);
  AN2 AND2_4143(g17317,g1079,g13124);
  AN2 AND2_4144(g22128,g6629,g19277);
  AN2 AND2_4145(g33352,g32237,g20712);
  AN4 AND4_253(I31207,g32754,g32755,g32756,g32757);
  AN2 AND2_4146(g16636,g5929,g14768);
  AN2 AND2_4147(g18629,g3680,g17226);
  AN2 AND2_4148(g25142,g4717,g22885);
  AN2 AND2_4149(g18451,g2295,g15224);
  AN2 AND2_4150(g26347,g262,g24850);
  AN2 AND2_4151(g18472,g2413,g15224);
  AN2 AND2_4152(g32414,g4944,g30999);
  AN2 AND2_4153(g29188,g27163,g12762);
  AN2 AND2_4154(g33418,g32372,g21425);
  AN2 AND2_4155(g33822,g33385,g20157);
  AN2 AND2_4156(g18220,g1002,g16100);
  AN2 AND2_4157(g26253,g2327,g25435);
  AN2 AND2_4158(g30006,g29032,g9259);
  AN2 AND2_4159(g31266,g30129,g27742);
  AN2 AND2_4160(g31170,g19128,g29814);
  AN2 AND2_4161(g21452,g16119,g13624);
  AN2 AND2_4162(g18628,g15095,g17226);
  AN2 AND2_4163(g27427,g26400,g17575);
  AN2 AND2_4164(g34475,g27450,g34327);
  AN2 AND2_4165(g17057,g446,g13173);
  AN2 AND2_4166(g24140,g17663,g21654);
  AN2 AND2_4167(g22299,g19999,g21024);
  AN2 AND2_4168(g29686,g2246,g29057);
  AN2 AND2_4169(g24997,g22929,g10419);
  AN2 AND2_4170(g18246,g1199,g16431);
  AN2 AND2_4171(g21912,g5052,g21468);
  AN2 AND2_4172(g29383,g28138,g19412);
  AN2 AND2_4173(g30222,g28701,g23894);
  AN2 AND2_4174(g34863,g16540,g34833);
  AN2 AND2_4175(g28133,g27367,g23108);
  AN2 AND2_4176(g22298,g19997,g21012);
  AN4 AND4_254(g26236,g25357,g6856,g7586,g7558);
  AN2 AND2_4177(g28229,g27345,g17213);
  AN2 AND2_4178(g19487,g499,g16680);
  AN2 AND2_4179(g29938,g23552,g28889);
  AN2 AND2_4180(g26351,g239,g24869);
  AN2 AND2_4181(g28228,g27126,g19636);
  AN2 AND2_4182(g25130,g23358,g20600);
  AN2 AND2_4183(g26821,g24821,g13103);
  AN2 AND2_4184(g27661,g26576,g15568);
  AN4 AND4_255(I31241,g30825,g31838,g32803,g32804);
  AN2 AND2_4185(g27547,g26549,g17759);
  AN2 AND2_4186(g18591,g2965,g16349);
  AN2 AND2_4187(g31194,g19128,g29814);
  AN2 AND2_4188(g31167,g10080,g30076);
  AN2 AND2_4189(g18776,g5813,g18065);
  AN2 AND2_4190(g18785,g5849,g18065);
  AN2 AND2_4191(g15083,g10362,g12983);
  AN2 AND2_4192(g21756,g3211,g20785);
  AN2 AND2_4193(g18147,g599,g17533);
  AN2 AND2_4194(g25165,g14062,g23570);
  AN2 AND2_4195(g30253,g28746,g23943);
  AN2 AND2_4196(g16484,g5244,g14755);
  AN2 AND2_4197(g18754,g5339,g15595);
  AN2 AND2_4198(g31524,g29897,g20593);
  AN3 AND3_234(g33524,g32918,I31316,I31317);
  AN2 AND2_4199(g18355,g1748,g17955);
  AN4 AND4_256(g26264,g24688,g8812,g8778,g10627);
  AN2 AND2_4200(g33836,g33096,g27020);
  AN2 AND2_4201(g21780,g3391,g20391);
  AN2 AND2_4202(g29875,g28403,g23337);
  AN2 AND2_4203(g32206,g30609,g25524);
  AN2 AND2_4204(g26516,g24968,g8876);
  AN2 AND2_4205(g13507,g7023,g12198);
  AN2 AND2_4206(g27481,g26400,g14630);
  AN2 AND2_4207(g30600,g30287,g18975);
  AN2 AND2_4208(g18825,g6736,g15680);
  AN2 AND2_4209(g18950,g11193,g16123);
  AN2 AND2_4210(g18370,g1874,g15171);
  AN2 AND2_4211(g31477,g29763,g23409);
  AN2 AND2_4212(g33401,g32349,g21381);
  AN3 AND3_235(g33477,g32577,I31081,I31082);
  AN2 AND2_4213(g20162,g8737,g16750);
  AN2 AND2_4214(g30236,g28724,g23916);
  AN2 AND2_4215(g14148,g884,g10632);
  AN2 AND2_4216(g29837,g28369,g20144);
  AN2 AND2_4217(g14097,g878,g10632);
  AN2 AND2_4218(g21820,g3712,g20453);
  AN2 AND2_4219(g11163,g6727,g10224);
  AN3 AND3_236(I24067,g3731,g3736,g8553);
  AN2 AND2_4220(g9906,g996,g1157);
  AN2 AND2_4221(g18151,g617,g17533);
  AN2 AND2_4222(g31118,g29490,g22906);
  AN2 AND2_4223(g18172,g15058,g17328);
  AN2 AND2_4224(g28627,g27543,g20574);
  AN2 AND2_4225(g32114,g31624,g29927);
  AN4 AND4_257(g28959,g17401,g25194,g26424,g27440);
  AN2 AND2_4226(g30175,g28629,g23813);
  AN2 AND2_4227(g32082,g4917,g30673);
  AN2 AND2_4228(g33864,g33274,g20524);
  AN2 AND2_4229(g27127,g25997,g16582);
  AN2 AND2_4230(g21846,g3897,g21070);
  AN2 AND2_4231(g28112,g27352,g26162);
  AN2 AND2_4232(g32107,g31624,g29912);
  AN2 AND2_4233(g15653,g3119,g13530);
  AN2 AND2_4234(g24629,g6163,g23699);
  AN2 AND2_4235(g23396,g20051,g20229);
  AN2 AND2_4236(g18367,g1783,g17955);
  AN2 AND2_4237(g18394,g1862,g15171);
  AN2 AND2_4238(g31313,g30160,g27907);
  AN2 AND2_4239(g24451,g3476,g23112);
  AN2 AND2_4240(g21731,g3029,g20330);
  AN2 AND2_4241(g24220,g255,g22594);
  AN2 AND2_4242(g20628,g1046,g15789);
  AN2 AND2_4243(g27490,g26576,g17651);
  AN2 AND2_4244(g13541,g7069,g12308);
  AN2 AND2_4245(g30264,g28774,g23963);
  AN2 AND2_4246(g34063,g33806,g23121);
  AN2 AND2_4247(g13473,g9797,g11841);
  AN2 AND2_4248(g30137,g28594,g21181);
  AN2 AND2_4249(g19601,g16198,g11149);
  AN2 AND2_4250(g24628,g5835,g23666);
  AN2 AND2_4251(g32345,g2138,g31672);
  AN2 AND2_4252(g34137,g33928,g23802);
  AN2 AND2_4253(g31285,g30134,g27800);
  AN2 AND2_4254(g34516,g34289,g19492);
  AN2 AND2_4255(g27376,g26549,g17481);
  AN2 AND2_4256(g27385,g26400,g17497);
  AN3 AND3_237(g33704,g33176,g10710,g22319);
  AN2 AND2_4257(g29617,g2024,g28987);
  AN2 AND2_4258(g31305,g29741,g23354);
  AN4 AND4_258(I24695,g24050,g24051,g24052,g24053);
  AN3 AND3_238(I24018,g8155,g8390,g3396);
  AN2 AND2_4259(g27103,g25997,g16509);
  AN2 AND2_4260(g33305,g31935,g17811);
  AN2 AND2_4261(g22831,g19441,g19629);
  AN2 AND2_4262(g23691,g14731,g20993);
  AN2 AND2_4263(g26542,g13102,g24376);
  AN2 AND2_4264(g34873,g34830,g20046);
  AN2 AND2_4265(g26021,g9568,g25035);
  AN2 AND2_4266(g18420,g1996,g15373);
  AN2 AND2_4267(g15852,g13820,g13223);
  AN2 AND2_4268(g27095,g25997,g16473);
  AN2 AND2_4269(g18319,g1600,g17873);
  AN2 AND2_4270(g33809,g33432,g30184);
  AN2 AND2_4271(g33900,g33316,g20913);
  AN3 AND3_239(g33466,g32498,I31026,I31027);
  AN2 AND2_4272(g16184,g9285,g14183);
  AN2 AND2_4273(g16805,g7187,g12972);
  AN2 AND2_4274(g21405,g13377,g15811);
  AN2 AND2_4275(g16674,g6637,g15014);
  AN3 AND3_240(g29201,g24081,I27503,I27504);
  AN2 AND2_4276(g32141,g31639,g29963);
  AN2 AND2_4277(g22316,g2837,g20270);
  AN2 AND2_4278(g18318,g1604,g17873);
  AN2 AND2_4279(g18446,g2279,g18008);
  AN2 AND2_4280(g33808,g33109,g22161);
  AN2 AND2_4281(g24785,g7051,g23645);
  AN2 AND2_4282(g18227,g1052,g16129);
  AN3 AND3_241(g7777,g723,g822,g817);
  AN2 AND2_4283(g27181,g26026,g16655);
  AN2 AND2_4284(g30209,g28682,g23876);
  AN3 AND3_242(g22498,g7753,g7717,g21334);
  AN2 AND2_4285(g33101,g32398,g18976);
  AN2 AND2_4286(g19791,g14253,g17189);
  AN2 AND2_4287(g24754,g19604,g23027);
  AN2 AND2_4288(g29595,g28475,g11833);
  AN2 AND2_4289(g29494,g9073,g28479);
  AN2 AND2_4290(g30208,g28681,g23875);
  AN2 AND2_4291(g16732,g5555,g14882);
  AN2 AND2_4292(g21929,g5176,g18997);
  AN2 AND2_4293(g32263,g31631,g30306);
  AN2 AND2_4294(g18540,g2775,g15277);
  AN2 AND2_4295(g10896,g1205,g8654);
  AN2 AND2_4296(g22056,g6133,g21611);
  AN2 AND2_4297(g26274,g2130,g25210);
  AN2 AND2_4298(g29623,g28496,g11563);
  AN2 AND2_4299(g32332,g31325,g23558);
  AN4 AND4_259(I31206,g31710,g31832,g32752,g32753);
  AN2 AND2_4300(g21928,g5170,g18997);
  AN2 AND2_4301(g22080,g6275,g19210);
  AN2 AND2_4302(g25063,g13078,g22325);
  AN3 AND3_243(g24858,g3361,g23223,I24030);
  AN2 AND2_4303(g29782,g28328,g23245);
  AN2 AND2_4304(g18203,g911,g15938);
  AN2 AND2_4305(g26122,g24557,g19762);
  AN2 AND2_4306(g16761,g7170,g12947);
  AN2 AND2_4307(g29984,g2567,g28877);
  AN2 AND2_4308(g34542,g34332,g20089);
  AN3 AND3_244(g22432,g9354,g7717,g21187);
  AN2 AND2_4309(g12931,g392,g11048);
  AN2 AND2_4310(g29352,g4950,g28410);
  AN2 AND2_4311(g25873,g24854,g16197);
  AN2 AND2_4312(g30614,g20154,g29814);
  AN3 AND3_245(I24597,g5736,g5742,g9875);
  AN4 AND4_260(I31082,g32573,g32574,g32575,g32576);
  AN2 AND2_4313(g18281,g1373,g16136);
  AN2 AND2_4314(g27520,g26519,g17714);
  AN2 AND2_4315(g21787,g15091,g20391);
  AN2 AND2_4316(g15115,g2946,g14454);
  AN4 AND4_261(I31107,g32610,g32611,g32612,g32613);
  AN3 AND3_246(g22342,g9354,g9285,g21287);
  AN2 AND2_4317(g18301,g1532,g16489);
  AN2 AND2_4318(g30607,g30291,g18989);
  AN2 AND2_4319(g32049,g10902,g30735);
  AN4 AND4_262(I24689,g20841,g24040,g24041,g24042);
  AN2 AND2_4320(g26292,g2689,g25228);
  AN2 AND2_4321(g33693,g33145,g13594);
  AN2 AND2_4322(g18377,g1894,g15171);
  AN2 AND2_4323(g19556,g11932,g16809);
  AN2 AND2_4324(g30073,g1379,g28194);
  AN2 AND2_4325(g22145,g14555,g18832);
  AN2 AND2_4326(g18120,g457,g17015);
  AN2 AND2_4327(g26153,g24565,g19780);
  AN2 AND2_4328(g18739,g5008,g16826);
  AN2 AND2_4329(g21302,g956,g15731);
  AN2 AND2_4330(g22031,g5917,g19147);
  AN2 AND2_4331(g27546,g26549,g17758);
  AN2 AND2_4332(g30274,g28815,g23983);
  AN2 AND2_4333(g31166,g1816,g30074);
  AN2 AND2_4334(g34073,g8948,g33823);
  AN2 AND2_4335(g10925,g7858,g956);
  AN2 AND2_4336(g16207,g9839,g14204);
  AN2 AND2_4337(g27211,g25997,g16716);
  AN2 AND2_4338(g32048,g31498,g13869);
  AN4 AND4_263(g16539,g11547,g6782,g6789,I17741);
  AN2 AND2_4339(g21743,g3100,g20330);
  AN2 AND2_4340(g21827,g3759,g20453);
  AN2 AND2_4341(g11029,g5782,g9103);
  AN2 AND2_4342(g17753,g13281,g13175);
  AN2 AND2_4343(g18146,g595,g17533);
  AN2 AND2_4344(g18738,g15142,g16826);
  AN2 AND2_4345(g13029,g8359,g11030);
  AN2 AND2_4346(g15745,g686,g13223);
  AN2 AND2_4347(g18645,g15100,g17271);
  AN2 AND2_4348(g30122,g28578,g21054);
  AN2 AND2_4349(g24420,g23997,g18980);
  AN2 AND2_4350(g24319,g4561,g22228);
  AN2 AND2_4351(g29853,g1862,g29081);
  AN2 AND2_4352(g16538,g6255,g15005);
  AN2 AND2_4353(g17145,g7469,g13249);
  AN2 AND2_4354(g26635,g25321,g20617);
  AN2 AND2_4355(g11028,g9730,g5428);
  AN2 AND2_4356(g18699,g4760,g16816);
  AN2 AND2_4357(g34565,g34374,g17471);
  AN2 AND2_4358(g15813,g3247,g14069);
  AN2 AND2_4359(g31485,g29776,g23421);
  AN2 AND2_4360(g29589,g2575,g28977);
  AN2 AND2_4361(g33892,g33312,g20701);
  AN2 AND2_4362(g18290,g1467,g16449);
  AN2 AND2_4363(g17199,g2236,g13034);
  AN2 AND2_4364(g24318,g4555,g22228);
  AN3 AND3_247(g33476,g32570,I31076,I31077);
  AN3 AND3_248(g33485,g32635,I31121,I31122);
  AN2 AND2_4365(g21769,g3247,g20785);
  AN2 AND2_4366(g30034,g29077,g10541);
  AN2 AND2_4367(g22843,g9429,g20272);
  AN2 AND2_4368(g24227,g890,g22594);
  AN2 AND2_4369(g18698,g15131,g16777);
  AN4 AND4_264(I31141,g31376,g31820,g32659,g32660);
  AN3 AND3_249(g25453,g5406,g23789,I24576);
  AN2 AND2_4370(g29588,g2311,g28942);
  AN2 AND2_4371(g29524,g2004,g28864);
  AN2 AND2_4372(g29836,g28425,g26841);
  AN2 AND2_4373(g21768,g3243,g20785);
  AN2 AND2_4374(g21803,g3538,g20924);
  AN2 AND2_4375(g28245,g11367,g27975);
  AN2 AND2_4376(g15805,g3243,g14041);
  AN2 AND2_4377(g28626,g27542,g20573);
  AN2 AND2_4378(g30153,g28610,g23768);
  AN2 AND2_4379(g28299,g9716,g27670);
  AN4 AND4_265(g27700,g22342,g25182,g26424,g26148);
  AN2 AND2_4380(g22132,g6645,g19277);
  AN2 AND2_4381(g29477,g14090,g28441);
  AN2 AND2_4382(g32273,g31255,g20446);
  AN2 AND2_4383(g32106,g31601,g29911);
  AN2 AND2_4384(g18427,g2181,g18008);
  AN2 AND2_4385(g14681,g4392,g10476);
  AN2 AND2_4386(g19740,g2783,g15907);
  AN2 AND2_4387(g20203,g6195,g17789);
  AN3 AND3_250(g33907,g23088,g33219,g9104);
  AN2 AND2_4388(g18366,g1854,g17955);
  AN4 AND4_266(I31332,g32935,g32936,g32937,g32938);
  AN2 AND2_4389(g21881,g4064,g19801);
  AN2 AND2_4390(g27658,g22491,g25786);
  AN2 AND2_4391(g18632,g3698,g17226);
  AN2 AND2_4392(g25905,g24879,g16311);
  AN2 AND2_4393(g17365,g7650,g13036);
  AN2 AND2_4394(g22161,g13202,g19071);
  AN2 AND2_4395(g33074,g32387,g18830);
  AN2 AND2_4396(g34136,g33850,g23293);
  AN2 AND2_4397(g33239,g32117,g19902);
  AN2 AND2_4398(g25530,g23750,g21414);
  AN2 AND2_4399(g27339,g26400,g17308);
  AN2 AND2_4400(g29749,g28295,g23214);
  AN2 AND2_4401(g29616,g1974,g29085);
  AN3 AND3_251(g7511,g2145,g2138,g2130);
  AN2 AND2_4402(g26711,g25446,g20713);
  AN2 AND2_4403(g31238,g29583,g20053);
  AN2 AND2_4404(g32234,g31601,g30292);
  AN2 AND2_4405(g25122,g23374,g20592);
  AN2 AND2_4406(g18403,g2028,g15373);
  AN2 AND2_4407(g18547,g121,g15277);
  AN2 AND2_4408(g25565,g13013,g22660);
  AN2 AND2_4409(g24301,g6961,g22228);
  AN2 AND2_4410(g28232,g27732,g23586);
  AN2 AND2_4411(g20739,g16259,g4674);
  AN2 AND2_4412(g13491,g6999,g12160);
  AN2 AND2_4413(g22087,g6303,g19210);
  AN2 AND2_4414(g30164,g28618,g23787);
  AN2 AND2_4415(g31941,g1283,g30825);
  AN2 AND2_4416(g33941,g33380,g21560);
  AN2 AND2_4417(g18226,g15064,g16129);
  AN2 AND2_4418(g21890,g4125,g19801);
  AN2 AND2_4419(g13604,g4495,g10487);
  AN2 AND2_4420(g31519,g29864,g23490);
  AN2 AND2_4421(g18715,g4871,g15915);
  AN2 AND2_4422(g27968,g25958,g19614);
  AN2 AND2_4423(g28697,g27581,g20669);
  AN2 AND2_4424(g31185,g10114,g30087);
  AN2 AND2_4425(g18481,g2461,g15426);
  AN3 AND3_252(g33519,g32881,I31291,I31292);
  AN2 AND2_4426(g29809,g28362,g23274);
  AN3 AND3_253(g33675,g33164,g10727,g22332);
  AN2 AND2_4427(g24645,g22639,g19709);
  AN2 AND2_4428(g28261,g27878,g23695);
  AN2 AND2_4429(g26606,g1018,g24510);
  AN4 AND4_267(g28880,g21434,g26424,g25438,g27494);
  AN2 AND2_4430(g18551,g2811,g15277);
  AN2 AND2_4431(g22043,g5965,g19147);
  AN2 AND2_4432(g26303,g2685,g25439);
  AN2 AND2_4433(g31518,g20041,g29970);
  AN2 AND2_4434(g31154,g19128,g29814);
  AN2 AND2_4435(g18572,g2864,g16349);
  AN3 AND3_254(g33518,g32874,I31286,I31287);
  AN2 AND2_4436(g29808,g28361,g23273);
  AN2 AND2_4437(g21710,g287,g20283);
  AN4 AND4_268(I31221,g31327,g31835,g32773,g32774);
  AN2 AND2_4438(g24290,g4430,g22550);
  AN4 AND4_269(g29036,g27163,g12762,g20875,I27381);
  AN2 AND2_4439(g27411,g26549,g17528);
  AN2 AND2_4440(g34474,g20083,g34326);
  AN2 AND2_4441(g24698,g22664,g19761);
  AN2 AND2_4442(g21779,g3385,g20391);
  AN2 AND2_4443(g26750,g24514,g24474);
  AN2 AND2_4444(g12527,g8680,g667);
  AN2 AND2_4445(g23779,g1105,g19355);
  AN2 AND2_4446(g18127,g499,g16971);
  AN2 AND2_4447(g22069,g6227,g19210);
  AN2 AND2_4448(g25408,g22682,g9772);
  AN2 AND2_4449(g30109,g28562,g20912);
  AN2 AND2_4450(g26381,g4456,g25548);
  AN2 AND2_4451(g34109,g33918,g23708);
  AN2 AND2_4452(g29642,g27954,g28669);
  AN2 AND2_4453(g33883,g33294,g20589);
  AN2 AND2_4454(g21778,g3355,g20391);
  AN2 AND2_4455(g22068,g6219,g19210);
  AN2 AND2_4456(g26091,g1691,g25082);
  AN2 AND2_4457(g18490,g2504,g15426);
  AN2 AND2_4458(g30108,g28561,g20910);
  AN2 AND2_4459(g32163,g3502,g31170);
  AN2 AND2_4460(g32012,g8297,g31233);
  AN3 AND3_255(g34108,g22957,g9104,g33766);
  AN2 AND2_4461(g24427,g4961,g22919);
  AN2 AND2_4462(g21786,g3436,g20391);
  AN2 AND2_4463(g27503,g26488,g14668);
  AN3 AND3_256(I24054,g8443,g8075,g3747);
  AN2 AND2_4464(g30283,g28851,g23993);
  AN4 AND4_270(I31106,g30825,g31814,g32608,g32609);
  AN2 AND2_4465(g18784,g15155,g18065);
  AN2 AND2_4466(g18376,g1913,g15171);
  AN2 AND2_4467(g18385,g1959,g15171);
  AN2 AND2_4468(g29733,g2675,g29157);
  AN2 AND2_4469(g18297,g1478,g16449);
  AN2 AND2_4470(g17810,g1495,g13246);
  AN2 AND2_4471(g18103,g401,g17015);
  AN2 AND2_4472(g10626,g4057,g7927);
  AN2 AND2_4473(g34492,g34272,g33430);
  AN2 AND2_4474(g13633,g4567,g10509);
  AN2 AND2_4475(g25164,g16883,g23569);
  AN2 AND2_4476(g21945,g5248,g18997);
  AN2 AND2_4477(g28499,g27982,g17762);
  AN2 AND2_4478(g18354,g1792,g17955);
  AN2 AND2_4479(g29874,g28402,g23336);
  AN4 AND4_271(g27714,g22384,g25195,g26424,g26171);
  AN2 AND2_4480(g21826,g3742,g20453);
  AN2 AND2_4481(g21999,g5723,g21562);
  AN2 AND2_4482(g26390,g4423,g25554);
  AN2 AND2_4483(g31501,g2047,g29310);
  AN2 AND2_4484(g18824,g6732,g15680);
  AN2 AND2_4485(g27315,g12022,g26709);
  AN3 AND3_257(g33501,g32751,I31201,I31202);
  AN2 AND2_4486(g29630,g28212,g19781);
  AN2 AND2_4487(g24403,g4894,g22858);
  AN2 AND2_4488(g29693,g28207,g10233);
  AN2 AND2_4489(g30982,g8895,g29933);
  AN2 AND2_4490(g34750,g34673,g19542);
  AN2 AND2_4491(g16759,g5587,g14761);
  AN2 AND2_4492(g18181,g772,g17328);
  AN2 AND2_4493(g21998,g5712,g21562);
  AN2 AND2_4494(g18671,g4628,g15758);
  AN2 AND2_4495(g34381,g34166,g20594);
  AN2 AND2_4496(g23998,g19631,g10971);
  AN3 AND3_258(g33728,g22626,g10851,g33187);
  AN2 AND2_4497(g27202,g25997,g13876);
  AN2 AND2_4498(g19568,g1467,g15959);
  AN2 AND2_4499(g30091,g28127,g20716);
  AN2 AND2_4500(g32325,g31316,g23538);
  AN2 AND2_4501(g29665,g2375,g28696);
  AN2 AND2_4502(g16758,g5220,g14758);
  AN3 AND3_259(g34091,g22957,g9104,g33761);
  AN2 AND2_4503(g24226,g446,g22594);
  AN2 AND2_4504(g13832,g8880,g10612);
  AN2 AND2_4505(g28722,g27955,g20738);
  AN4 AND4_272(g28924,g17317,g25183,g26424,g27416);
  AN2 AND2_4506(g30174,g28628,g23812);
  AN4 AND4_273(g29008,g27163,g12730,g20739,I27364);
  AN2 AND2_4507(g12979,g424,g11048);
  AN2 AND2_4508(g24551,g17148,g23331);
  AN2 AND2_4509(g24572,g5462,g23393);
  AN2 AND2_4510(g33349,g32233,g20699);
  AN2 AND2_4511(g25108,g23345,g20576);
  AN2 AND2_4512(g21932,g5204,g18997);
  AN2 AND2_4513(g32121,g31616,g29942);
  AN2 AND2_4514(g18426,g2177,g18008);
  AN2 AND2_4515(g33906,g33084,g22311);
  AN2 AND2_4516(g13247,g8964,g11316);
  AN2 AND2_4517(g29555,g29004,g22498);
  AN2 AND2_4518(g21513,g16196,g10882);
  AN2 AND2_4519(g18190,g822,g17821);
  AN2 AND2_4520(g22010,g5787,g21562);
  AN2 AND2_4521(g23513,g19430,g13007);
  AN2 AND2_4522(g34390,g34172,g21069);
  AN2 AND2_4523(g10856,g4269,g8967);
  AN2 AND2_4524(g11045,g5787,g9883);
  AN2 AND2_4525(g15882,g3554,g13986);
  AN2 AND2_4526(g27384,g26400,g17496);
  AN2 AND2_4527(g29570,g2763,g28598);
  AN2 AND2_4528(g29712,g2643,g28726);
  AN4 AND4_274(I24694,g20982,g24047,g24048,g24049);
  AN2 AND2_4529(g33304,g32427,g31971);
  AN2 AND2_4530(g14261,g4507,g10738);
  AN2 AND2_4531(g18520,g2661,g15509);
  AN2 AND2_4532(g21961,g5424,g21514);
  AN2 AND2_4533(g22079,g6271,g19210);
  AN2 AND2_4534(g27094,g25997,g16472);
  AN2 AND2_4535(g30192,g28649,g23847);
  AN2 AND2_4536(g31566,g19050,g29814);
  AN2 AND2_4537(g13324,g854,g11326);
  AN2 AND2_4538(g29907,g2629,g29177);
  AN2 AND2_4539(g32291,g31268,g20527);
  AN2 AND2_4540(g16804,g5905,g14813);
  AN2 AND2_4541(g21404,g16069,g13569);
  AN2 AND2_4542(g28199,g27479,g16684);
  AN2 AND2_4543(g22078,g6267,g19210);
  AN2 AND2_4544(g23404,g20063,g20247);
  AN2 AND2_4545(g32173,g160,g31134);
  AN2 AND2_4546(g18546,g2795,g15277);
  AN2 AND2_4547(g25982,g2351,g25008);
  AN4 AND4_275(I31012,g32473,g32474,g32475,g32476);
  AN2 AND2_4548(g18211,g15062,g15979);
  AN2 AND2_4549(g21717,g15051,g21037);
  AN2 AND2_4550(g28198,g26649,g27492);
  AN2 AND2_4551(g24297,g4455,g22550);
  AN2 AND2_4552(g22086,g6299,g19210);
  AN2 AND2_4553(g25091,g12830,g23492);
  AN2 AND2_4554(g20095,g8873,g16632);
  AN3 AND3_260(I24619,g6423,g6428,g10014);
  AN2 AND2_4555(g29567,g2357,g28593);
  AN2 AND2_4556(g29594,g28529,g14192);
  AN3 AND3_261(g12735,g7121,g3873,g3881);
  AN2 AND2_4557(g31139,g12221,g30036);
  AN2 AND2_4558(g28528,g27187,g12730);
  AN2 AND2_4559(g28330,g27238,g19786);
  AN2 AND2_4560(g26252,g2283,g25309);
  AN2 AND2_4561(g11032,g9354,g7717);
  AN2 AND2_4562(g34483,g34406,g18938);
  AN2 AND2_4563(g18497,g2541,g15426);
  AN2 AND2_4564(g32029,g31318,g16482);
  AN2 AND2_4565(g24671,g5481,g23630);
  AN2 AND2_4566(g14831,g1152,g10909);
  AN2 AND2_4567(g22125,g6617,g19277);
  AN3 AND3_262(g29382,g26424,g22763,g28172);
  AN2 AND2_4568(g27526,g26576,g17721);
  AN2 AND2_4569(g34862,g16540,g34830);
  AN2 AND2_4570(g29519,g2295,g28840);
  AN2 AND2_4571(g32028,g30569,g29339);
  AN2 AND2_4572(g19578,g16183,g11130);
  AN2 AND2_4573(g33415,g32368,g21422);
  AN2 AND2_4574(g22158,g13698,g19609);
  AN2 AND2_4575(g14316,g2370,g11920);
  AN2 AND2_4576(g33333,g32218,g20612);
  AN2 AND2_4577(g18700,g15132,g16816);
  AN4 AND4_276(g17817,g11547,g6782,g11640,I18819);
  AN2 AND2_4578(g18126,g15054,g16971);
  AN2 AND2_4579(g18659,g4366,g17183);
  AN2 AND2_4580(g18625,g15092,g17062);
  AN2 AND2_4581(g18987,g182,g16162);
  AN2 AND2_4582(g29518,g28906,g22384);
  AN2 AND2_4583(g18250,g6821,g16897);
  AN2 AND2_4584(g24931,g23153,g20178);
  AN2 AND2_4585(g15114,g4239,g14454);
  AN2 AND2_4586(g25192,g20276,g23648);
  AN2 AND2_4587(g26847,g2873,g24525);
  AN2 AND2_4588(g34948,g16540,g34935);
  AN2 AND2_4589(g18658,g15121,g17183);
  AN2 AND2_4590(g27457,g26519,g17606);
  AN2 AND2_4591(g26397,g19475,g25563);
  AN2 AND2_4592(g15082,g2697,g12983);
  AN2 AND2_4593(g23387,g16506,g20211);
  AN2 AND2_4594(g31963,g30731,g18895);
  AN2 AND2_4595(g29637,g2533,g29134);
  AN2 AND2_4596(g22680,g19530,g7781);
  AN2 AND2_4597(g34702,g34537,g20208);
  AN2 AND2_4598(g15107,g4258,g14454);
  AN2 AND2_4599(g23148,g19128,g9104);
  AN2 AND2_4600(g34757,g34682,g19635);
  AN2 AND2_4601(g17783,g7851,g13110);
  AN2 AND2_4602(g25522,g6888,g22544);
  AN4 AND4_277(I31121,g30614,g31817,g32629,g32630);
  AN2 AND2_4603(g24190,g329,g22722);
  AN2 AND2_4604(g18339,g1714,g17873);
  AN2 AND2_4605(g18943,g269,g16099);
  AN2 AND2_4606(g29883,g2465,g29152);
  AN2 AND2_4607(g18296,g1495,g16449);
  AN2 AND2_4608(g21811,g3582,g20924);
  AN2 AND2_4609(g28225,g27770,g23400);
  AN2 AND2_4610(g23104,g661,g20248);
  AN2 AND2_4611(g23811,g4087,g19364);
  AN2 AND2_4612(g23646,g16959,g20737);
  AN2 AND2_4613(g18644,g15098,g17125);
  AN4 AND4_278(g28471,g27187,g12762,g21024,I26960);
  AN2 AND2_4614(g16221,g5791,g14231);
  AN2 AND2_4615(g18338,g1710,g17873);
  AN2 AND2_4616(g30564,g21358,g29385);
  AN2 AND2_4617(g9967,g1178,g1157);
  AN2 AND2_4618(g28258,g27182,g19687);
  AN2 AND2_4619(g21971,g5417,g21514);
  AN2 AND2_4620(g34564,g34373,g17466);
  AN2 AND2_4621(g15849,g3538,g14136);
  AN2 AND2_4622(g31484,g29775,g23418);
  AN2 AND2_4623(g24546,g22447,g19523);
  AN3 AND3_263(g33484,g32628,I31116,I31117);
  AN2 AND2_4624(g16613,g5925,g14732);
  AN4 AND4_279(I31291,g31021,g31847,g32875,g32876);
  AN2 AND2_4625(g15848,g3259,g13892);
  AN2 AND2_4626(g19275,g7823,g16044);
  AN2 AND2_4627(g31554,g19050,g29814);
  AN2 AND2_4628(g30673,g20175,g29814);
  AN2 AND2_4629(g27256,g25937,g19698);
  AN2 AND2_4630(g19746,g9816,g17147);
  AN2 AND2_4631(g28244,g27926,g26715);
  AN2 AND2_4632(g34183,g33695,g24385);
  AN2 AND2_4633(g18197,g854,g17821);
  AN2 AND2_4634(g22017,g5763,g21562);
  AN2 AND2_4635(g15652,g174,g13437);
  AN2 AND2_4636(g15804,g3223,g13889);
  AN2 AND2_4637(g34397,g7673,g34068);
  AN2 AND2_4638(g25949,g24701,g19559);
  AN2 AND2_4639(g27280,g9825,g26614);
  AN2 AND2_4640(g31312,g30136,g27858);
  AN2 AND2_4641(g29577,g2441,g28946);
  AN2 AND2_4642(g30062,g13129,g28174);
  AN2 AND2_4643(g27300,g12370,g26672);
  AN2 AND2_4644(g10736,g4040,g8751);
  AN3 AND3_264(g10887,g7812,g6565,g6573);
  AN2 AND2_4645(g31115,g29487,g22882);
  AN2 AND2_4646(g18411,g2093,g15373);
  AN2 AND2_4647(g25536,g23770,g21431);
  AN2 AND2_4648(g25040,g12738,g23443);
  AN4 AND4_280(g26213,g25357,g11724,g7586,g7558);
  AN2 AND2_4649(g34509,g34283,g19473);
  AN2 AND2_4650(g21850,g3893,g21070);
  AN2 AND2_4651(g28602,g27509,g20515);
  AN2 AND2_4652(g23412,g7297,g21510);
  AN2 AND2_4653(g28657,g27562,g20606);
  AN2 AND2_4654(g25904,g14001,g24791);
  AN3 AND3_265(g33921,g33187,g9104,g19200);
  AN2 AND2_4655(g19684,g2735,g17297);
  AN2 AND2_4656(g34508,g34282,g19472);
  AN2 AND2_4657(g10528,g1576,g9051);
  AN2 AND2_4658(g34872,g34827,g19954);
  AN3 AND3_266(I18740,g13156,g11450,g11498);
  AN2 AND2_4659(g24700,g645,g23512);
  AN4 AND4_281(g28970,g17405,g25196,g26424,g27445);
  AN2 AND2_4660(g24659,g5134,g23590);
  AN4 AND4_282(g14528,g12459,g12306,g12245,I16646);
  AN2 AND2_4661(g26205,g2098,g25492);
  AN2 AND2_4662(g23229,g18994,g4521);
  AN4 AND4_283(g16234,g6772,g6782,g11640,I17575);
  AN2 AND2_4663(g29349,g4760,g28391);
  AN2 AND2_4664(g22309,g1478,g19751);
  AN2 AND2_4665(g20658,g1389,g15800);
  AN2 AND2_4666(g18503,g2563,g15509);
  AN2 AND2_4667(g22023,g5881,g19147);
  AN2 AND2_4668(g26311,g2527,g25400);
  AN2 AND2_4669(g24658,g22645,g19732);
  AN3 AND3_267(I24015,g8334,g7975,g3045);
  AN3 AND3_268(g10869,g7766,g5873,g5881);
  AN2 AND2_4670(g22308,g1135,g19738);
  AN2 AND2_4671(g28171,g27016,g19385);
  AN2 AND2_4672(g33798,g33227,g20058);
  AN2 AND2_4673(g21716,g301,g20283);
  AN2 AND2_4674(g30213,g28688,g23880);
  AN2 AND2_4675(g24296,g4382,g22550);
  AN2 AND2_4676(g18581,g2912,g16349);
  AN2 AND2_4677(g18714,g4864,g15915);
  AN2 AND2_4678(g26051,g24896,g14169);
  AN2 AND2_4679(g18450,g2299,g15224);
  AN2 AND2_4680(g31184,g1950,g30085);
  AN2 AND2_4681(g34213,g33766,g22689);
  AN2 AND2_4682(g18315,g1548,g16931);
  AN2 AND2_4683(g33805,g33232,g20079);
  AN3 AND3_269(g33674,g33164,g10710,g22319);
  AN2 AND2_4684(g24644,g11714,g22903);
  AN2 AND2_4685(g29622,g2579,g29001);
  AN2 AND2_4686(g29566,g2307,g28907);
  AN2 AND2_4687(g18707,g15134,g16782);
  AN2 AND2_4688(g18819,g6541,g15483);
  AN2 AND2_4689(g18910,g16227,g16075);
  AN2 AND2_4690(g18202,g907,g15938);
  AN2 AND2_4691(g30047,g29109,g9407);
  AN2 AND2_4692(g18257,g1205,g16897);
  AN2 AND2_4693(g26780,g4098,g24437);
  AN2 AND2_4694(g30205,g28671,g23869);
  AN2 AND2_4695(g32191,g27593,g31376);
  AN2 AND2_4696(g18818,g15165,g15483);
  AN2 AND2_4697(g18496,g2537,g15426);
  AN2 AND2_4698(g34205,g33729,g24541);
  AN2 AND2_4699(g31934,g31670,g18827);
  AN2 AND2_4700(g18111,g174,g17015);
  AN2 AND2_4701(g21959,g5413,g21514);
  AN2 AND2_4702(g21925,g5073,g21468);
  AN2 AND2_4703(g26350,g13087,g25517);
  AN2 AND2_4704(g25872,g3119,g24655);
  AN2 AND2_4705(g28919,g27663,g21295);
  AN2 AND2_4706(g14708,g74,g12369);
  AN3 AND3_270(I18762,g13156,g6767,g11498);
  AN4 AND4_284(g28458,g27187,g12730,g20887,I26948);
  AN2 AND2_4707(g24197,g347,g22722);
  AN3 AND3_271(g24855,g3050,g23534,I24027);
  AN3 AND3_272(g27660,g24688,g26424,g22763);
  AN2 AND2_4708(g16163,g14254,g14179);
  AN2 AND2_4709(g22752,g15792,g19612);
  AN2 AND2_4710(g15613,g3490,g13555);
  AN2 AND2_4711(g18590,g2917,g16349);
  AN2 AND2_4712(g21958,g5396,g21514);
  AN2 AND2_4713(g21378,g7887,g16090);
  AN2 AND2_4714(g23050,g655,g20248);
  AN4 AND4_285(g28010,g23032,g26223,g26424,g25535);
  AN2 AND2_4715(g23958,g9104,g19200);
  AN2 AND2_4716(g24411,g4584,g22161);
  AN2 AND2_4717(g30051,g28513,g20604);
  AN2 AND2_4718(g26846,g37,g24524);
  AN2 AND2_4719(g18741,g15143,g17384);
  AN2 AND2_4720(g34072,g33839,g24872);
  AN2 AND2_4721(g23386,g20034,g20207);
  AN2 AND2_4722(g30592,g30270,g18929);
  AN2 AND2_4723(g18384,g1945,g15171);
  AN2 AND2_4724(g29636,g2403,g29097);
  AN2 AND2_4725(g21742,g3050,g20330);
  AN2 AND2_4726(g17752,g7841,g13174);
  AN2 AND2_4727(g27480,g26400,g17638);
  AN2 AND2_4728(g34756,g34680,g19618);
  AN2 AND2_4729(g23742,g19128,g9104);
  AN2 AND2_4730(g28599,g27027,g8922);
  AN2 AND2_4731(g21944,g5244,g18997);
  AN2 AND2_4732(g33400,g32347,g21380);
  AN2 AND2_4733(g29852,g1772,g29080);
  AN2 AND2_4734(g17643,g9681,g14599);
  AN2 AND2_4735(g15812,g3227,g13915);
  AN4 AND4_286(g13319,g4076,g8812,g10658,g8757);
  AN2 AND2_4736(g27314,g12436,g26702);
  AN2 AND2_4737(g24503,g22225,g19409);
  AN2 AND2_4738(g27287,g26545,g23011);
  AN2 AND2_4739(g32045,g31491,g16187);
  AN4 AND4_287(I24685,g24036,g24037,g24038,g24039);
  AN2 AND2_4740(g33329,g32210,g20585);
  AN2 AND2_4741(g31207,g30252,g20739);
  AN2 AND2_4742(g18150,g604,g17533);
  AN2 AND2_4743(g10657,g8451,g4064);
  AN2 AND2_4744(g18801,g15160,g15348);
  AN2 AND2_4745(g18735,g4983,g16826);
  AN2 AND2_4746(g25574,I24709,I24710);
  AN2 AND2_4747(g27085,g25835,g22494);
  AN2 AND2_4748(g32324,g31315,g23537);
  AN2 AND2_4749(g29664,g2273,g29060);
  AN2 AND2_4750(g33328,g32209,g20584);
  AN2 AND2_4751(g21802,g3562,g20924);
  AN2 AND2_4752(g22489,g12954,g19386);
  AN2 AND2_4753(g21857,g3933,g21070);
  AN2 AND2_4754(g23802,g9104,g19050);
  AN2 AND2_4755(g16535,g5595,g14848);
  AN2 AND2_4756(g20581,g10801,g15571);
  AN2 AND2_4757(g10970,g854,g9582);
  AN2 AND2_4758(g23857,g19626,g7908);
  AN2 AND2_4759(g13059,g6900,g11303);
  AN2 AND2_4760(g13025,g8431,g11026);
  AN2 AND2_4761(g30152,g28609,g23767);
  AN2 AND2_4762(g24581,g5124,g23590);
  AN2 AND2_4763(g24714,g6173,g23699);
  AN2 AND2_4764(g32098,g4732,g30614);
  AN2 AND2_4765(g24450,g3129,g23067);
  AN2 AND2_4766(g21730,g3025,g20330);
  AN2 AND2_4767(g24315,g4521,g22228);
  AN2 AND2_4768(g21793,g3412,g20391);
  AN2 AND2_4769(g32272,g31639,g30310);
  AN2 AND2_4770(g22525,g13006,g19411);
  AN2 AND2_4771(g28159,g8553,g27317);
  AN4 AND4_288(I31262,g32833,g32834,g32835,g32836);
  AN2 AND2_4772(g10878,g7858,g1135);
  AN2 AND2_4773(g18196,g703,g17821);
  AN2 AND2_4774(g22016,g5747,g21562);
  AN2 AND2_4775(g28125,g27381,g26209);
  AN2 AND2_4776(g15795,g3566,g14130);
  AN2 AND2_4777(g18695,g4737,g16053);
  AN2 AND2_4778(g28532,g27394,g20265);
  AN2 AND2_4779(g34396,g34194,g21337);
  AN3 AND3_273(I18568,g13156,g11450,g11498);
  AN2 AND2_4780(g24707,g13295,g22997);
  AN2 AND2_4781(g30731,g11374,g29361);
  AN2 AND2_4782(g29576,g2177,g28903);
  AN2 AND2_4783(g29585,g1756,g28920);
  AN2 AND2_4784(g21765,g3231,g20785);
  AN3 AND3_274(g28158,g26424,g22763,g27037);
  AN4 AND4_289(I27523,g20857,g24111,g24112,g24113);
  AN2 AND2_4785(g18526,g2555,g15509);
  AN2 AND2_4786(g27269,g25943,g19734);
  AN2 AND2_4787(g29554,g28997,g22472);
  AN2 AND2_4788(g23690,g14726,g20978);
  AN2 AND2_4789(g19372,g686,g16289);
  AN2 AND2_4790(g26020,g9559,g25034);
  AN2 AND2_4791(g33241,g32173,g23128);
  AN2 AND2_4792(g34413,g34094,g22670);
  AN2 AND2_4793(g17424,g1426,g13176);
  AN2 AND2_4794(g11044,g5343,g10124);
  AN4 AND4_290(I31191,g30735,g31829,g32731,g32732);
  AN2 AND2_4795(g27341,g10203,g26788);
  AN2 AND2_4796(g10967,g7880,g1448);
  AN2 AND2_4797(g29609,g28482,g11861);
  AN2 AND2_4798(g27268,g25942,g19733);
  AN2 AND2_4799(g32032,g31373,g16515);
  AN2 AND2_4800(g25780,g25532,g25527);
  AN2 AND2_4801(g15507,g10970,g13305);
  AN2 AND2_4802(g32140,g31609,g29961);
  AN2 AND2_4803(g28144,g4608,g27020);
  AN2 AND2_4804(g18402,g2047,g15373);
  AN2 AND2_4805(g18457,g2319,g15224);
  AN2 AND2_4806(g24590,g6154,g23413);
  AN2 AND2_4807(g29608,g28568,g11385);
  AN2 AND2_4808(g27180,g26026,g16654);
  AN2 AND2_4809(g19516,g7824,g16097);
  AN2 AND2_4810(g20094,g8872,g16631);
  AN2 AND2_4811(g27335,g12087,g26776);
  AN3 AND3_275(g33683,g33149,g10727,g22332);
  AN2 AND2_4812(g13738,g8880,g10572);
  AN2 AND2_4813(g25152,g23383,g20626);
  AN2 AND2_4814(g22042,g5961,g19147);
  AN2 AND2_4815(g26302,g2393,g25349);
  AN2 AND2_4816(g26357,g22547,g25525);
  AN2 AND2_4817(g29799,g28271,g10233);
  AN2 AND2_4818(g30583,g19666,g29355);
  AN2 AND2_4819(g16760,g5559,g14764);
  AN2 AND2_4820(g27667,g26361,g20601);
  AN4 AND4_291(I31247,g32812,g32813,g32814,g32815);
  AN2 AND2_4821(g18706,g4785,g16782);
  AN2 AND2_4822(g18597,g2975,g16349);
  AN2 AND2_4823(g27965,g25834,g13117);
  AN2 AND2_4824(g13290,g3897,g11534);
  AN2 AND2_4825(g29798,g28348,g23260);
  AN2 AND2_4826(g22124,g6613,g19277);
  AN2 AND2_4827(g27131,g26055,g16588);
  AN2 AND2_4828(g30046,g29108,g10564);
  AN2 AND2_4829(g18256,g1242,g16897);
  AN2 AND2_4830(g29973,g28981,g9206);
  AN2 AND2_4831(g18689,g15129,g16752);
  AN2 AND2_4832(g31991,g4912,g30673);
  AN3 AND3_276(g33515,g32853,I31271,I31272);
  AN2 AND2_4833(g33882,g33293,g20587);
  AN2 AND2_4834(g18280,g1367,g16136);
  AN2 AND2_4835(g29805,g28357,g23270);
  AN2 AND2_4836(g33414,g32367,g21421);
  AN2 AND2_4837(g22686,g19335,g19577);
  AN2 AND2_4838(g22939,g9708,g21062);
  AN2 AND2_4839(g18688,g4704,g16752);
  AN2 AND2_4840(g18624,g3490,g17062);
  AN2 AND2_4841(g32162,g31002,g23014);
  AN2 AND2_4842(g18300,g1306,g16489);
  AN2 AND2_4843(g24196,g333,g22722);
  AN2 AND2_4844(g33407,g32357,g21406);
  AN2 AND2_4845(g34113,g33734,g19744);
  AN2 AND2_4846(g27502,g26488,g17677);
  AN4 AND4_292(I31251,g31710,g31840,g32817,g32818);
  AN2 AND2_4847(g11427,g5706,g7158);
  AN2 AND2_4848(g22030,g5909,g19147);
  AN4 AND4_293(I31272,g32849,g32850,g32851,g32852);
  AN2 AND2_4849(g22938,g19782,g19739);
  AN2 AND2_4850(g27557,g26549,g17774);
  AN2 AND2_4851(g22093,g6423,g18833);
  AN2 AND2_4852(g23533,g19436,g13015);
  AN2 AND2_4853(g11366,g5016,g10338);
  AN3 AND3_277(g27210,g26218,g8373,g2476);
  AN2 AND2_4854(g21298,g7697,g15825);
  AN2 AND2_4855(g29732,g2514,g29131);
  AN2 AND2_4856(g28289,g27734,g26575);
  AN2 AND2_4857(g21775,g3372,g20391);
  AN3 AND3_278(I16671,g10185,g12461,g12415);
  AN2 AND2_4858(g13632,g10232,g12228);
  AN2 AND2_4859(g18157,g15057,g17433);
  AN2 AND2_4860(g23775,g14872,g21267);
  AN2 AND2_4861(g22065,g6203,g19210);
  AN3 AND3_279(g34105,g33778,g9104,g18957);
  AN3 AND3_280(g28224,g27163,g22763,g27064);
  AN2 AND2_4862(g34743,g8951,g34703);
  AN3 AND3_281(I17585,g14988,g11450,g11498);
  AN2 AND2_4863(g28571,g27458,g20435);
  AN2 AND2_4864(g24402,g4749,g22857);
  AN2 AND2_4865(g29761,g28310,g23228);
  AN4 AND4_294(I31032,g32501,g32502,g32503,g32504);
  AN2 AND2_4866(g18231,g1105,g16326);
  AN2 AND2_4867(g21737,g3068,g20330);
  AN2 AND2_4868(g32246,g31246,g20326);
  AN4 AND4_295(g27469,g8046,g26314,g518,g9077);
  AN2 AND2_4869(g22219,g19953,g20887);
  AN2 AND2_4870(g25928,g25022,g23436);
  AN2 AND2_4871(g8583,g2917,g2912);
  AN2 AND2_4872(g27286,g6856,g26634);
  AN2 AND2_4873(g33441,g32251,g29722);
  AN2 AND2_4874(g31206,g30260,g23890);
  AN2 AND2_4875(g10656,g3782,g7952);
  AN4 AND4_296(g27039,g7738,g5527,g5535,g26223);
  AN2 AND2_4876(g22218,g19951,g20875);
  AN2 AND2_4877(g28495,g27012,g12465);
  AN2 AND2_4878(g32071,g27236,g31070);
  AN4 AND4_297(I31061,g30825,g31806,g32543,g32544);
  AN2 AND2_4879(g21856,g3929,g21070);
  AN3 AND3_282(g10823,g7704,g5180,g5188);
  AN2 AND2_4880(g14295,g1811,g11894);
  AN2 AND2_4881(g21995,g5611,g19074);
  AN2 AND2_4882(g31759,g21291,g29385);
  AN2 AND2_4883(g23856,g4116,g19483);
  AN2 AND2_4884(g14680,g12024,g12053);
  AN2 AND2_4885(g33759,g33123,g22847);
  AN3 AND3_283(g33725,g22626,g10851,g33176);
  AN2 AND2_4886(g24001,g19651,g10951);
  AN2 AND2_4887(g21880,g4135,g19801);
  AN2 AND2_4888(g29329,g7995,g28353);
  AN2 AND2_4889(g25113,g23346,g20577);
  AN2 AND2_4890(g18511,g2599,g15509);
  AN3 AND3_284(g29207,g24131,I27533,I27534);
  AN2 AND2_4891(g25787,g24792,g20887);
  AN2 AND2_4892(g32147,g31616,g29980);
  AN2 AND2_4893(g18763,g5481,g17929);
  AN2 AND2_4894(g31758,g30115,g23945);
  AN2 AND2_4895(g33114,g22139,g31945);
  AN2 AND2_4896(g24706,g15910,g22996);
  AN2 AND2_4897(g26249,g1858,g25300);
  AN2 AND2_4898(g33758,g33133,g20269);
  AN2 AND2_4899(g22160,g8005,g19795);
  AN2 AND2_4900(g27601,g26766,g26737);
  AN2 AND2_4901(g33082,g32389,g18877);
  AN2 AND2_4902(g21512,g16225,g10881);
  AN3 AND3_285(g29328,g28553,g6928,g3990);
  AN2 AND2_4903(g27677,g13021,g25888);
  AN2 AND2_4904(g25357,g23810,g23786);
  AN2 AND2_4905(g29538,g2563,g28914);
  AN2 AND2_4906(g11127,g6479,g10022);
  AN2 AND2_4907(g24923,g23129,g20167);
  AN2 AND2_4908(g25105,g13973,g23505);
  AN2 AND2_4909(g10966,g9226,g7948);
  AN2 AND2_4910(g31744,g30092,g23902);
  AN2 AND2_4911(g24688,g22681,g22663);
  AN2 AND2_4912(g26204,g1720,g25275);
  AN2 AND2_4913(g24624,g16524,g22867);
  AN2 AND2_4914(g24300,g15123,g22228);
  AN3 AND3_286(I24579,g5731,g5736,g9875);
  AN2 AND2_4915(g26779,g24497,g23620);
  AN2 AND2_4916(g33345,g32229,g20671);
  AN2 AND2_4917(g32151,g31639,g29996);
  AN2 AND2_4918(g32172,g2767,g31608);
  AN4 AND4_298(I31162,g32689,g32690,g32691,g32692);
  AN2 AND2_4919(g31940,g943,g30735);
  AN2 AND2_4920(g18456,g2338,g15224);
  AN2 AND2_4921(g33849,g33262,g20387);
  AN2 AND2_4922(g30027,g29104,g12550);
  AN2 AND2_4923(g33399,g32346,g21379);
  AN2 AND2_4924(g21831,g3782,g20453);
  AN2 AND2_4925(g26778,g25501,g20923);
  AN2 AND2_4926(g34662,g34576,g18931);
  AN2 AND2_4927(g16845,g6593,g15011);
  AN2 AND2_4928(g11956,g2070,g7411);
  AN2 AND2_4929(g18480,g2437,g15426);
  OR2 OR2_0(g32367,g29880,g31309);
  OR2 OR2_1(g34890,g34863,g21674);
  OR2 OR2_2(g28668,g27411,g16617);
  OR2 OR2_3(g34249,g34110,g21702);
  OR2 OR2_4(g13095,g11374,g1287);
  OR2 OR2_5(g30482,g30230,g21978);
  OR2 OR2_6(g24231,g22589,g18201);
  OR2 OR2_7(g13888,g2941,g11691);
  OR2 OR2_8(g26945,g26379,g24283);
  OR2 OR2_9(g30552,g30283,g22123);
  OR2 OR2_10(g34003,g33866,g18452);
  OR2 OR2_11(g23989,g20581,g17179);
  OR2 OR2_12(g29235,g28110,g18260);
  OR2 OR2_13(g28525,g27284,g26176);
  OR2 OR2_14(g34204,g33832,g33833);
  OR4 OR4_0(I28566,g29201,g29202,g29203,g28035);
  OR2 OR2_15(g14309,g10320,g11048);
  OR4 OR4_1(I30330,g29385,g31376,g30735,g30825);
  OR2 OR2_16(g24854,g21453,g24002);
  OR2 OR2_17(g30081,g28454,g11366);
  OR2 OR2_18(g32227,g31146,g29648);
  OR2 OR2_19(g33962,g33822,g18123);
  OR2 OR2_20(g19575,g15693,g13042);
  OR2 OR2_21(g27556,g26097,g24687);
  OR2 OR2_22(g25662,g24656,g21787);
  OR2 OR2_23(g28544,g27300,g26229);
  OR2 OR2_24(g30356,g30096,g18365);
  OR2 OR2_25(g27580,g26159,g24749);
  OR2 OR2_26(g34647,g34558,g18820);
  OR2 OR2_27(g26932,g26684,g18549);
  OR4 OR4_2(I31859,g33501,g33502,g33503,g33504);
  OR2 OR2_28(g33049,g31966,g21929);
  OR2 OR2_29(g30380,g30161,g18492);
  OR2 OR2_30(g34826,g34742,g34685);
  OR3 OR3_0(g16926,g14061,g11804,g11780);
  OR3 OR3_1(I25736,g12,g22150,g20277);
  OR4 OR4_3(I31858,g33497,g33498,g33499,g33500);
  OR2 OR2_31(g33048,g31960,g21928);
  OR2 OR2_32(g7684,g4072,g4176);
  OR2 OR2_33(g25710,g25031,g21961);
  OR2 OR2_34(g28610,g27347,g16484);
  OR2 OR2_35(g26897,g26611,g18176);
  OR2 OR2_36(g34090,g33676,g33680);
  OR2 OR2_37(g26961,g26280,g24306);
  OR2 OR2_38(g28705,g27460,g16672);
  OR2 OR2_39(g28042,g24148,g26879);
  OR2 OR2_40(g30672,g13737,g29752);
  OR2 OR2_41(g34233,g32455,g33951);
  OR2 OR2_42(g13211,g11294,g7567);
  OR2 OR2_43(g33004,g32246,g18431);
  OR2 OR2_44(g31221,g29494,g28204);
  OR3 OR3_2(g23198,g20214,g20199,I22298);
  OR4 OR4_4(I31844,g33474,g33475,g33476,g33477);
  OR2 OR2_45(g27179,g25816,g24409);
  OR2 OR2_46(g28188,g22535,g27108);
  OR2 OR2_47(g33613,g33248,g18649);
  OR2 OR2_48(g34331,g27121,g34072);
  OR2 OR2_49(g30513,g30200,g22034);
  OR2 OR2_50(g30449,g29845,g21858);
  OR2 OR2_51(g33947,g32438,g33457);
  OR2 OR2_52(g34449,g34279,g18662);
  OR2 OR2_53(g25647,g24725,g21740);
  OR2 OR2_54(g24243,g22992,g18254);
  OR2 OR2_55(g33273,g32122,g29553);
  OR2 OR2_56(g28030,g24018,g26874);
  OR2 OR2_57(g33605,g33352,g18521);
  OR2 OR2_58(g25945,g24427,g22307);
  OR2 OR2_59(g28093,g27981,g21951);
  OR2 OR2_60(g30448,g29809,g21857);
  OR2 OR2_61(g34897,g34861,g21682);
  OR2 OR2_62(g34448,g34365,g18553);
  OR2 OR2_63(g30505,g30168,g22026);
  OR2 OR2_64(g29114,g27646,g26602);
  OR2 OR2_65(g30404,g29758,g21763);
  OR2 OR2_66(g28065,g27299,g21792);
  OR2 OR2_67(g27800,g17321,g26703);
  OR2 OR2_68(g24269,g23131,g18613);
  OR2 OR2_69(g34404,g34182,g25102);
  OR3 OR3_3(g33951,g33469,I31838,I31839);
  OR2 OR2_70(g33972,g33941,g18335);
  OR2 OR2_71(g24341,g23564,g18771);
  OR2 OR2_72(g33033,g32333,g21843);
  OR2 OR2_73(g24268,g23025,g18612);
  OR2 OR2_74(g25651,g24680,g21744);
  OR2 OR2_75(g25672,g24647,g21829);
  OR2 OR2_76(g33234,g32039,g32043);
  OR2 OR2_77(g34026,g33715,g18682);
  OR2 OR2_78(g32427,g8928,g30583);
  OR2 OR2_79(g13296,g10626,g10657);
  OR2 OR2_80(g23087,g19487,g15852);
  OR2 OR2_81(g29849,g26049,g28273);
  OR2 OR2_82(g13969,g11448,g8913);
  OR2 OR2_83(g26343,g1514,g24609);
  OR2 OR2_84(g19522,g17057,g14180);
  OR2 OR2_85(g29848,g28260,g26077);
  OR2 OR2_86(g24335,g22165,g18678);
  OR2 OR2_87(g26971,g26325,g24333);
  OR2 OR2_88(g34723,g34710,g18139);
  OR2 OR2_89(g30433,g29899,g21817);
  OR2 OR2_90(g34149,g33760,g19674);
  OR2 OR2_91(g30387,g30151,g18524);
  OR2 OR2_92(g24965,g22667,g23825);
  OR2 OR2_93(g32226,g31145,g29645);
  OR2 OR2_94(g29263,g28239,g18617);
  OR2 OR2_95(g34620,g34529,g18582);
  OR2 OR2_96(g34148,g33758,g19656);
  OR2 OR2_97(g25717,g25106,g21968);
  OR2 OR2_98(g27543,g26085,g24670);
  OR2 OR2_99(g30104,g28478,g11427);
  OR2 OR2_100(g33012,g32274,g18483);
  OR2 OR2_101(g19949,g17671,g14681);
  OR2 OR2_102(g30343,g29344,g18278);
  OR2 OR2_103(g34646,g34557,g18803);
  OR2 OR2_104(g24557,g22308,g19207);
  OR2 OR2_105(g24210,g22900,g18125);
  OR2 OR2_106(g27569,g26124,g24721);
  OR2 OR2_107(g34971,g34869,g34962);
  OR2 OR2_108(g33541,g33101,g18223);
  OR2 OR2_109(g31473,g26180,g29666);
  OR2 OR2_110(g28075,g27083,g21877);
  OR2 OR2_111(g30369,g30066,g18439);
  OR2 OR2_112(g24443,g23917,g21378);
  OR2 OR2_113(g19904,g17636,g14654);
  OR2 OR2_114(g23171,g19536,g15903);
  OR2 OR2_115(g24279,g23218,g15105);
  OR2 OR2_116(g26896,g26341,g18171);
  OR2 OR2_117(g34369,g26279,g34136);
  OR2 OR2_118(g28595,g27335,g26290);
  OR2 OR2_119(g14030,g11037,g11046);
  OR2 OR2_120(g30368,g30098,g18435);
  OR2 OR2_121(g24278,g23201,g18648);
  OR2 OR2_122(g25723,g25033,g22006);
  OR2 OR2_123(g28623,g27361,g16520);
  OR2 OR2_124(g34368,g26274,g34135);
  OR2 OR2_125(g33788,g33122,g32041);
  OR2 OR2_126(g31325,g29625,g29639);
  OR2 OR2_127(g32385,g31480,g29938);
  OR2 OR2_128(g31920,g31493,g22045);
  OR2 OR2_129(g32980,g32254,g18198);
  OR2 OR2_130(g30412,g29885,g21771);
  OR2 OR2_131(g33535,g33233,g21711);
  OR2 OR2_132(g24468,g10925,g22400);
  OR2 OR2_133(g32354,g29854,g31285);
  OR2 OR2_134(g34850,g34841,g18185);
  OR2 OR2_135(g34412,g34187,g25143);
  OR2 OR2_136(g28419,g27221,g15884);
  OR2 OR2_137(g27974,g26544,g25063);
  OR2 OR2_138(g33946,g32434,g33456);
  OR2 OR2_139(g25646,g24706,g21739);
  OR2 OR2_140(g28418,g27220,g15882);
  OR2 OR2_141(g20187,g16202,g13491);
  OR2 OR2_142(g26959,g26381,g24299);
  OR2 OR2_143(g26925,g25939,g18301);
  OR2 OR2_144(g34011,g33884,g18479);
  OR2 OR2_145(g26958,g26395,g24297);
  OR2 OR2_146(g29273,g28269,g18639);
  OR2 OR2_147(g31291,g29581,g29593);
  OR4 OR4_5(g17570,g14419,g14397,g11999,I18495);
  OR2 OR2_148(g33291,g32154,g13477);
  OR2 OR2_149(g26386,g24719,g23023);
  OR3 OR3_4(g32426,g26105,g26131,g30613);
  OR2 OR2_150(g28194,g22540,g27122);
  OR2 OR2_151(g28589,g27331,g26285);
  OR2 OR2_152(g26944,g26130,g18658);
  OR2 OR2_153(g20169,g16184,g13460);
  OR2 OR2_154(g27579,g26157,g24748);
  OR2 OR2_155(g29234,g28415,g18239);
  OR2 OR2_156(g30379,g30089,g18491);
  OR2 OR2_157(g34627,g34534,g18644);
  OR2 OR2_158(g27578,g26155,g24747);
  OR4 OR4_6(g17594,g14450,g14420,g12025,I18543);
  OR2 OR2_159(g28401,g27212,g15871);
  OR2 OR2_160(g31760,g30007,g30027);
  OR2 OR2_161(g34379,g26312,g34143);
  OR2 OR2_162(g33029,g32332,g21798);
  OR2 OR2_163(g32211,g31124,g29603);
  OR2 OR2_164(g30378,g30125,g18487);
  OR2 OR2_165(g21901,g21251,g15115);
  OR2 OR2_166(g20217,g16221,g13523);
  OR2 OR2_167(g33028,g32325,g21797);
  OR2 OR2_168(g30386,g30139,g18523);
  OR2 OR2_169(g24363,g7831,g22138);
  OR2 OR2_170(g26793,g24478,g7520);
  OR2 OR2_171(g28118,g27821,g26815);
  OR3 OR3_5(g13526,g209,g10685,g301);
  OR2 OR2_172(g24478,g11003,g22450);
  OR2 OR2_173(g34603,g34561,g15075);
  OR2 OR2_174(g25716,g25088,g21967);
  OR2 OR2_175(g28749,g27523,g16764);
  OR2 OR2_176(g26690,g10776,g24433);
  OR2 OR2_177(g25582,g21662,g24152);
  OR2 OR2_178(g28748,g27522,g16763);
  OR2 OR2_179(g28704,g27459,g16671);
  OR2 OR2_180(g24580,g22340,g13096);
  OR2 OR2_181(g31927,g31500,g22091);
  OR2 OR2_182(g30429,g29844,g21813);
  OR2 OR2_183(g28305,g27103,g15793);
  OR2 OR2_184(g28053,g27393,g18168);
  OR2 OR2_185(g32987,g32311,g18323);
  OR2 OR2_186(g32250,g30598,g29351);
  OR2 OR2_187(g34802,g34757,g18589);
  OR2 OR2_188(g25627,g24503,g18247);
  OR2 OR2_189(g30428,g29807,g21812);
  OR2 OR2_190(g34730,g34658,g18271);
  OR2 OR2_191(g34793,g34744,g18570);
  OR4 OR4_7(I26643,g27073,g27058,g27045,g27040);
  OR2 OR2_192(g13077,g11330,g943);
  OR3 OR3_6(I18492,g14538,g14513,g14446);
  OR2 OR2_193(g28101,g27691,g22062);
  OR2 OR2_194(g33240,g32052,g32068);
  OR2 OR2_195(g13597,g9247,g11149);
  OR2 OR2_196(g28560,g27311,g26249);
  OR2 OR2_197(g31903,g31374,g21911);
  OR2 OR2_198(g30549,g30215,g22120);
  OR2 OR2_199(g25603,g24698,g18114);
  OR2 OR2_200(g25742,g25093,g22057);
  OR2 OR2_201(g31755,g29991,g30008);
  OR2 OR2_202(g33604,g33345,g18520);
  OR2 OR2_203(g30548,g30204,g22119);
  OR2 OR2_204(g10589,g7223,g7201);
  OR2 OR2_205(g29325,g28813,g27820);
  OR2 OR2_206(g13300,g10656,g10676);
  OR2 OR2_207(g31770,g30034,g30047);
  OR2 OR2_208(g30504,g30253,g22025);
  OR2 OR2_209(g28064,g27298,g21781);
  OR2 OR2_210(g33563,g33361,g18383);
  OR2 OR2_211(g33981,g33856,g18371);
  OR2 OR2_212(g25681,g24710,g18636);
  OR2 OR2_213(g28733,g27507,g16735);
  OR2 OR2_214(g26299,g24551,g22665);
  OR3 OR3_7(g30317,g29208,I28566,I28567);
  OR2 OR2_215(g25730,g25107,g22013);
  OR2 OR2_216(g22304,g21347,g17693);
  OR2 OR2_217(g14119,g10776,g8703);
  OR2 OR2_218(g31767,g30031,g30043);
  OR2 OR2_219(g33794,g33126,g32053);
  OR2 OR2_220(g34002,g33857,g18451);
  OR2 OR2_221(g33262,g32112,g29528);
  OR2 OR2_222(g31899,g31470,g21907);
  OR2 OR2_223(g34057,g33911,g33915);
  OR2 OR2_224(g28665,g27409,g16614);
  OR2 OR2_225(g30128,g28495,g11497);
  OR2 OR2_226(g33990,g33882,g18399);
  OR2 OR2_227(g24334,g23991,g18676);
  OR2 OR2_228(g25690,g24864,g21889);
  OR2 OR2_229(g26737,g24460,g10720);
  OR2 OR2_230(g29291,g28660,g18767);
  OR2 OR2_231(g31898,g31707,g21906);
  OR2 OR2_232(g34626,g34533,g18627);
  OR2 OR2_233(g30533,g30203,g22079);
  OR2 OR2_234(g22653,g18993,g15654);
  OR2 OR2_235(g30298,g28245,g27251);
  OR3 OR3_8(g23687,g21384,g21363,I22830);
  OR2 OR2_236(g26880,g26610,g24186);
  OR2 OR2_237(g24216,g23416,g18197);
  OR2 OR2_238(g23374,g19767,g13514);
  OR2 OR2_239(g32202,g31069,g13410);
  OR2 OR2_240(g22636,g18943,g15611);
  OR2 OR2_241(g26512,g24786,g23130);
  OR2 OR2_242(g32257,g31184,g29708);
  OR2 OR2_243(g13660,g8183,g12527);
  OR2 OR2_244(g32979,g32181,g18177);
  OR2 OR2_245(g29506,g28148,g25880);
  OR2 OR2_246(g34232,g33451,g33944);
  OR2 OR2_247(g32978,g32197,g18145);
  OR2 OR2_248(g28074,g27119,g21876);
  OR2 OR2_249(g33573,g33343,g18415);
  OR2 OR2_250(g31247,g29513,g13324);
  OR2 OR2_251(g28594,g27334,g26289);
  OR2 OR2_252(g31926,g31765,g22090);
  OR2 OR2_253(g32986,g31996,g18280);
  OR2 OR2_254(g27253,g24661,g26052);
  OR2 OR2_255(g33389,g32272,g29964);
  OR2 OR2_256(g33045,g32206,g24328);
  OR2 OR2_257(g22664,g19139,g15694);
  OR2 OR2_258(g34856,g34811,g34743);
  OR2 OR2_259(g25626,g24499,g18235);
  OR2 OR2_260(g33612,g33247,g18633);
  OR2 OR2_261(g34261,g34074,g18688);
  OR2 OR2_262(g34880,g34867,g18153);
  OR2 OR2_263(g8921,I12902,I12903);
  OR2 OR2_264(g30512,g30191,g22033);
  OR2 OR2_265(g33534,g33186,g21700);
  OR2 OR2_266(g27236,g24620,g25974);
  OR2 OR2_267(g32094,g30612,g29363);
  OR2 OR2_268(g31251,g25973,g29527);
  OR2 OR2_269(g22585,g20915,g21061);
  OR2 OR2_270(g33251,g32096,g29509);
  OR2 OR2_271(g24242,g22834,g18253);
  OR2 OR2_272(g33272,g32121,g29551);
  OR2 OR2_273(g28092,g27666,g21924);
  OR4 OR4_8(I30124,g31070,g31154,g30614,g30673);
  OR2 OR2_274(g28518,g27281,g26158);
  OR2 OR2_275(g21893,g20094,g18655);
  OR2 OR2_276(g29240,g28655,g18328);
  OR2 OR2_277(g26080,g19393,g24502);
  OR3 OR3_9(I12583,g1157,g1239,g990);
  OR2 OR2_278(g25737,g25045,g22052);
  OR2 OR2_279(g26924,g26153,g18291);
  OR2 OR2_280(g30445,g29772,g21854);
  OR2 OR2_281(g33032,g32326,g21842);
  OR2 OR2_282(g34445,g34382,g18548);
  OR2 OR2_283(g30499,g30261,g21995);
  OR2 OR2_284(g33997,g33871,g18427);
  OR2 OR2_285(g25697,g25086,g21916);
  OR4 OR4_9(g25856,g25518,g25510,g25488,g25462);
  OR2 OR2_286(g30498,g30251,g21994);
  OR2 OR2_287(g25261,g23348,g20193);
  OR2 OR2_288(g33061,g32334,g22050);
  OR2 OR2_289(g24265,g22316,g18560);
  OR2 OR2_290(g26342,g8407,g24591);
  OR2 OR2_291(g31766,g30029,g30042);
  OR2 OR2_292(g31871,g30596,g18279);
  OR2 OR2_293(g30611,g13671,g29743);
  OR2 OR2_294(g24841,g21420,g23998);
  OR2 OR2_295(g34611,g34508,g18565);
  OR2 OR2_296(g23255,g19655,g16122);
  OR2 OR2_297(g34722,g34707,g18137);
  OR2 OR2_298(g26887,g26542,g24193);
  OR2 OR2_299(g28729,g27502,g16732);
  OR2 OR2_300(g28577,g27326,g26272);
  OR2 OR2_301(g24510,g22488,g7567);
  OR2 OR2_302(g30432,g29888,g21816);
  OR2 OR2_303(g28728,g27501,g16730);
  OR2 OR2_304(g29262,g28327,g18608);
  OR2 OR2_305(g27542,g16190,g26094);
  OR2 OR2_306(g27453,g25976,g24606);
  OR2 OR2_307(g23383,g19756,g16222);
  OR2 OR2_308(g24578,g2882,g23825);
  OR2 OR2_309(g30461,g30219,g21932);
  OR2 OR2_310(g30342,g29330,g18261);
  OR2 OR2_311(g34461,g34291,g18681);
  OR2 OR2_312(g26365,g25504,g25141);
  OR3 OR3_10(I18452,g14514,g14448,g14418);
  OR2 OR2_313(g26960,g26258,g24304);
  OR2 OR2_314(g34031,g33735,g18705);
  OR2 OR2_315(g31472,g29642,g28352);
  OR2 OR2_316(g28083,g27249,g18689);
  OR2 OR2_317(g28348,g27139,g15823);
  OR2 OR2_318(g34199,g33820,g33828);
  OR2 OR2_319(g32280,g24790,g31225);
  OR2 OR2_320(g9984,g4300,g4242);
  OR2 OR2_321(g34887,g34865,g21670);
  OR2 OR2_322(g31911,g31784,g21969);
  OR2 OR2_323(g30529,g30212,g22075);
  OR2 OR2_324(g33628,g33071,g32450);
  OR2 OR2_325(g27274,g15779,g25915);
  OR2 OR2_326(g31246,g25965,g29518);
  OR2 OR2_327(g25611,g24931,g18128);
  OR2 OR2_328(g19356,g17784,g14874);
  OR2 OR2_329(g25722,g25530,g18768);
  OR2 OR2_330(g28622,g27360,g16519);
  OR2 OR2_331(g28566,g27316,g26254);
  OR2 OR2_332(g30528,g30202,g22074);
  OR2 OR2_333(g9483,g1008,g969);
  OR2 OR2_334(g30393,g29986,g21748);
  OR2 OR2_335(g27122,g22537,g25917);
  OR2 OR2_336(g34843,g33924,g34782);
  OR2 OR2_337(g34330,g34069,g33717);
  OR2 OR2_338(g30365,g30158,g18412);
  OR2 OR2_339(g24275,g23474,g18645);
  OR2 OR2_340(g29247,g28694,g18410);
  OR2 OR2_341(g31591,g29358,g29353);
  OR2 OR2_342(g31785,g30071,g30082);
  OR2 OR2_343(g33591,g33082,g18474);
  OR2 OR2_344(g24430,g23151,g8234);
  OR2 OR2_345(g24746,g22588,g19461);
  OR2 OR2_346(g32231,g30590,g29346);
  OR2 OR2_347(g25753,g25165,g22100);
  OR2 OR2_348(g31754,g29989,g30006);
  OR2 OR2_349(g28138,g27964,g27968);
  OR2 OR2_350(g24237,g22515,g18242);
  OR2 OR2_351(g33950,g32450,g33460);
  OR2 OR2_352(g29777,g28227,g28234);
  OR2 OR2_353(g24340,g24016,g18770);
  OR2 OR2_354(g25650,g24663,g21743);
  OR2 OR2_355(g25736,g25536,g18785);
  OR2 OR2_356(g29251,g28679,g18464);
  OR2 OR2_357(g29272,g28346,g18638);
  OR2 OR2_358(g28636,g27376,g16538);
  OR2 OR2_359(g19449,g15567,g12939);
  OR2 OR2_360(g28852,g27559,g16871);
  OR2 OR2_361(g34259,g34066,g18679);
  OR2 OR2_362(g30471,g30175,g21942);
  OR2 OR2_363(g33996,g33862,g18426);
  OR2 OR2_364(g34708,g33381,g34572);
  OR4 OR4_10(g26657,g24908,g24900,g24887,g24861);
  OR2 OR2_365(g25696,g25012,g21915);
  OR2 OR2_366(g26955,g26391,g24293);
  OR2 OR2_367(g34258,g34211,g18675);
  OR2 OR2_368(g24517,g22158,g18906);
  OR2 OR2_369(g26879,g25580,g25581);
  OR2 OR2_370(g26970,g26308,g24332);
  OR2 OR2_371(g25764,g25551,g18819);
  OR2 OR2_372(g28664,g27408,g16613);
  OR2 OR2_373(g26878,g25578,g25579);
  OR2 OR2_374(g16867,g13493,g11045);
  OR2 OR2_375(g25960,g24566,g24678);
  OR2 OR2_376(g34043,g33903,g33905);
  OR2 OR2_377(g26886,g26651,g24192);
  OR2 OR2_378(g25868,g25450,g23885);
  OR2 OR2_379(g28576,g27325,g26271);
  OR2 OR2_380(g31319,g29612,g28324);
  OR2 OR2_381(g27575,g26147,g24731);
  OR2 OR2_382(g26967,g26350,g24319);
  OR2 OR2_383(g33318,g31969,g32434);
  OR2 OR2_384(g34602,g34489,g18269);
  OR2 OR2_385(g25709,g25014,g21960);
  OR2 OR2_386(g30375,g30149,g18466);
  OR2 OR2_387(g34657,g33114,g34497);
  OR2 OR2_388(g28609,g27346,g16483);
  OR2 OR2_389(g33227,g32029,g32031);
  OR2 OR2_390(g9536,g1351,g1312);
  OR2 OR2_391(g33059,g31987,g22021);
  OR2 OR2_392(g33025,g32162,g21780);
  OR2 OR2_393(g25708,g25526,g18751);
  OR2 OR2_394(g34970,g34868,g34961);
  OR4 OR4_11(I29986,g31070,g31194,g30614,g30673);
  OR2 OR2_395(g23822,g20218,g16929);
  OR2 OR2_396(g33540,g33099,g18207);
  OR2 OR2_397(g27108,g22522,g25911);
  OR2 OR2_398(g33058,g31976,g22020);
  OR2 OR2_399(g30337,g29334,g18220);
  OR2 OR2_400(g32243,g31166,g29683);
  OR2 OR2_401(g26919,g25951,g18267);
  OR2 OR2_402(g28052,g27710,g18167);
  OR2 OR2_403(g27283,g25922,g25924);
  OR2 OR2_404(g26918,g25931,g18243);
  OR2 OR2_405(g28745,g27519,g16760);
  OR2 OR2_406(g15968,g13038,g10677);
  OR4 OR4_12(I31854,g33492,g33493,g33494,g33495);
  OR2 OR2_407(g33044,g32199,g24327);
  OR2 OR2_408(g34792,g34750,g18569);
  OR2 OR2_409(g32268,g24785,g31219);
  OR2 OR2_410(g23194,g19564,g19578);
  OR2 OR2_411(g33281,g32142,g29576);
  OR2 OR2_412(g31902,g31744,g21910);
  OR2 OR2_413(g30459,g29314,g21926);
  OR2 OR2_414(g30425,g29770,g21809);
  OR3 OR3_11(g33957,g33523,I31868,I31869);
  OR2 OR2_415(g24347,g23754,g18790);
  OR2 OR2_416(g34459,g34415,g18673);
  OR2 OR2_417(g25602,g24673,g18113);
  OR2 OR2_418(g12982,g12220,g9968);
  OR2 OR2_419(g25657,g24624,g21782);
  OR2 OR2_420(g24253,g22525,g18300);
  OR2 OR2_421(g25774,g25223,g12043);
  OR2 OR2_422(g29246,g28710,g18406);
  OR2 OR2_423(g30458,g30005,g24330);
  OR2 OR2_424(g34458,g34396,g18671);
  OR2 OR2_425(g33562,g33414,g18379);
  OR2 OR2_426(g34010,g33872,g18478);
  OR2 OR2_427(g24236,g22489,g18241);
  OR2 OR2_428(g25878,g25503,g23920);
  OR2 OR2_429(g28732,g27505,g16734);
  OR2 OR2_430(g33699,g32409,g33433);
  OR2 OR2_431(g32993,g32255,g18352);
  OR2 OR2_432(g30545,g30268,g22116);
  OR2 OR2_433(g30444,g29901,g21853);
  OR2 OR2_434(g29776,g28225,g22846);
  OR3 OR3_12(g24952,g21326,g21340,I24117);
  OR2 OR2_435(g24351,g23774,g18807);
  OR2 OR2_436(g33290,g32149,g29589);
  OR2 OR2_437(g26901,g26362,g24218);
  OR2 OR2_438(g34444,g34389,g18546);
  OR2 OR2_439(g24821,g21404,g23990);
  OR2 OR2_440(g29754,g28215,g28218);
  OR2 OR2_441(g34599,g34542,g18149);
  OR2 OR2_442(g32131,g24495,g30926);
  OR2 OR2_443(g20063,g15978,g13313);
  OR2 OR2_444(g34598,g34541,g18136);
  OR2 OR2_445(g15910,g13025,g10654);
  OR2 OR2_446(g24264,g22310,g18559);
  OR2 OR2_447(g23276,g19681,g16161);
  OR2 OR2_448(g27663,g26323,g24820);
  OR2 OR2_449(g28400,g27211,g15870);
  OR2 OR2_450(g32210,g31123,g29600);
  OR2 OR2_451(g21900,g20977,g15114);
  OR2 OR2_452(g16866,g13492,g11044);
  OR2 OR2_453(g28329,g27128,g15813);
  OR2 OR2_454(g30532,g30193,g22078);
  OR2 OR2_455(g32279,g31220,g31224);
  OR2 OR2_456(g34125,g33724,g33124);
  OR2 OR2_457(g22652,g18992,g15653);
  OR2 OR2_458(g13762,g499,g12527);
  OR2 OR2_459(g34977,g34873,g34966);
  OR2 OR2_460(g25010,g23267,g2932);
  OR2 OR2_461(g31895,g31505,g24296);
  OR2 OR2_462(g28328,g27127,g15812);
  OR2 OR2_463(g33547,g33349,g18331);
  OR2 OR2_464(g34158,g33784,g19740);
  OR2 OR2_465(g24209,g23415,g18122);
  OR2 OR2_466(g34783,g33110,g34667);
  OR2 OR2_467(g28538,g27294,g26206);
  OR2 OR2_468(g26966,g26345,g24318);
  OR2 OR2_469(g25545,g23551,g20658);
  OR2 OR2_470(g30561,g30284,g22132);
  OR2 OR2_471(g7673,g4153,g4172);
  OR2 OR2_472(g30353,g30095,g18355);
  OR2 OR2_473(g24208,g23404,g18121);
  OR2 OR2_474(g25599,g24914,g21721);
  OR2 OR2_475(g34353,g26088,g34114);
  OR2 OR2_476(g29319,g28812,g14453);
  OR2 OR2_477(g25598,g24904,g21720);
  OR2 OR2_478(g33551,g33446,g18342);
  OR2 OR2_479(g33572,g33339,g18414);
  OR2 OR2_480(g30336,g29324,g18203);
  OR2 OR2_481(g29227,g28456,g18169);
  OR2 OR2_482(g13543,g10543,g10565);
  OR4 OR4_13(I31839,g33465,g33466,g33467,g33468);
  OR4 OR4_14(I31838,g33461,g33462,g33463,g33464);
  OR2 OR2_483(g28100,g27690,g22051);
  OR2 OR2_484(g20905,g7216,g17264);
  OR2 OR2_485(g34631,g34562,g15118);
  OR2 OR2_486(g30364,g30086,g18411);
  OR2 OR2_487(g34017,g33880,g18504);
  OR2 OR2_488(g24274,g23187,g18631);
  OR2 OR2_489(g13242,g11336,g7601);
  OR3 OR3_13(g33956,g33514,I31863,I31864);
  OR2 OR2_490(g24346,g23725,g18789);
  OR2 OR2_491(g33297,g32157,g29621);
  OR2 OR2_492(g25656,g24945,g18609);
  OR2 OR2_493(g31889,g31118,g21822);
  OR2 OR2_494(g33980,g33843,g18370);
  OR2 OR2_495(g24565,g22309,g19275);
  OR2 OR2_496(g21892,g19788,g15104);
  OR2 OR2_497(g25680,g24794,g21839);
  OR3 OR3_14(g16876,g14028,g11773,g11755);
  OR2 OR2_498(g29281,g28541,g18743);
  OR2 OR2_499(g31888,g31067,g21821);
  OR2 OR2_500(g20034,g15902,g13299);
  OR2 OR2_501(g29301,g28686,g18797);
  OR2 OR2_502(g27509,g26023,g24640);
  OR2 OR2_503(g34289,g26847,g34218);
  OR2 OR2_504(g24641,g22151,g22159);
  OR2 OR2_505(g34023,g33796,g24320);
  OR2 OR2_506(g34288,g26846,g34217);
  OR2 OR2_507(g32217,g31129,g29616);
  OR2 OR2_508(g26954,g26380,g24292);
  OR3 OR3_15(I18449,g14512,g14445,g14415);
  OR2 OR2_509(g31931,g31494,g22095);
  OR2 OR2_510(g29290,g28569,g18764);
  OR2 OR2_511(g25631,g24554,g18275);
  OR2 OR2_512(g30495,g30222,g21991);
  OR2 OR2_513(g32223,g31142,g29637);
  OR2 OR2_514(g29366,g13738,g28439);
  OR2 OR2_515(g27574,g26145,g24730);
  OR2 OR2_516(g34976,g34872,g34965);
  OR2 OR2_517(g26392,g24745,g23050);
  OR2 OR2_518(g27205,g25833,g24421);
  OR2 OR2_519(g33546,g33402,g18327);
  OR2 OR2_520(g30374,g30078,g18465);
  OR2 OR2_521(g16076,g13081,g10736);
  OR2 OR2_522(g34374,g26294,g34139);
  OR4 OR4_15(I30728,g32345,g32350,g32056,g32018);
  OR2 OR2_523(g33024,g32324,g21752);
  OR2 OR2_524(g34643,g34554,g18752);
  OR2 OR2_525(g28435,g27234,g15967);
  OR2 OR2_526(g28082,g27369,g24315);
  OR2 OR2_527(g26893,g26753,g24199);
  OR2 OR2_528(g29226,g28455,g18159);
  OR2 OR2_529(g28744,g27518,g16759);
  OR2 OR2_530(g34260,g34113,g18680);
  OR2 OR2_531(g28345,g27137,g15821);
  OR2 OR2_532(g29481,g28117,g28125);
  OR2 OR2_533(g30392,g30091,g18558);
  OR2 OR2_534(g30489,g30250,g21985);
  OR2 OR2_535(g33625,g33373,g18809);
  OR2 OR2_536(g32373,g29894,g31321);
  OR2 OR2_537(g33987,g33847,g18396);
  OR2 OR2_538(g31250,g25972,g29526);
  OR2 OR2_539(g25687,g24729,g21882);
  OR2 OR2_540(g30559,g30269,g22130);
  OR2 OR2_541(g30525,g30266,g22071);
  OR2 OR2_542(g30488,g30197,g21984);
  OR2 OR2_543(g30424,g29760,g21808);
  OR2 OR2_544(g25752,g25079,g22099);
  OR2 OR2_545(g34016,g33867,g18503);
  OR2 OR2_546(g30558,g30258,g22129);
  OR2 OR2_547(g27152,g24393,g25817);
  OR2 OR2_548(g33296,g32156,g29617);
  OR2 OR2_549(g25643,g24602,g21736);
  OR2 OR2_550(g29490,g25832,g28136);
  OR2 OR2_551(g16839,g13473,g11035);
  OR2 OR2_552(g28332,g27130,g15815);
  OR2 OR2_553(g30544,g30257,g22115);
  OR2 OR2_554(g33969,g33864,g18321);
  OR2 OR2_555(g25669,g24657,g18624);
  OR2 OR2_556(g28135,g27959,g27963);
  OR2 OR2_557(g29297,g28683,g18784);
  OR2 OR2_558(g33060,g31992,g22022);
  OR2 OR2_559(g33968,g33855,g18320);
  OR2 OR2_560(g26939,g25907,g21884);
  OR2 OR2_561(g25668,g24646,g18623);
  OR3 OR3_16(g33197,g32342,I30745,I30746);
  OR2 OR2_562(g28361,g27153,g15839);
  OR2 OR2_563(g32216,g31128,g29615);
  OR2 OR2_564(g27405,g24572,g25968);
  OR2 OR2_565(g26938,g26186,g21883);
  OR2 OR2_566(g31870,g30607,g18262);
  OR3 OR3_17(I28147,g2946,g24561,g28220);
  OR2 OR2_567(g24840,g21419,g23996);
  OR2 OR2_568(g34610,g34507,g18564);
  OR2 OR2_569(g24390,g23779,g21285);
  OR2 OR2_570(g30189,g23401,g28543);
  OR2 OR2_571(g28049,g27684,g18164);
  OR2 OR2_572(g34255,g34120,g24302);
  OR2 OR2_573(g34189,g33801,g33808);
  OR2 OR2_574(g30270,g28624,g27664);
  OR2 OR2_575(g28048,g27362,g18163);
  OR2 OR2_576(g20522,g691,g16893);
  OR2 OR2_577(g26875,g21652,g25575);
  OR2 OR2_578(g32117,g24482,g30914);
  OR4 OR4_16(I23163,g20982,g21127,g21193,g21256);
  OR2 OR2_579(g31894,g30671,g21870);
  OR2 OR2_580(g31867,g31238,g18175);
  OR2 OR2_581(g30460,g30207,g21931);
  OR2 OR2_582(g30383,g30138,g18513);
  OR2 OR2_583(g34460,g34301,g18677);
  OR2 OR2_584(g30093,g28467,g11397);
  OR2 OR2_585(g34030,g33727,g18704);
  OR2 OR2_586(g25713,g25147,g21964);
  OR2 OR2_587(g28613,g27350,g26310);
  OR2 OR2_588(g33581,g33333,g18443);
  OR2 OR2_589(g33714,g32419,g33450);
  OR4 OR4_17(g29520,g28291,g28281,g28264,g28254);
  OR2 OR2_590(g34267,g34079,g18728);
  OR2 OR2_591(g34294,g26855,g34225);
  OR2 OR2_592(g31315,g29607,g29623);
  OR2 OR2_593(g33315,g29665,g32175);
  OR2 OR2_594(g31910,g31471,g21957);
  OR2 OR2_595(g13006,g12284,g10034);
  OR2 OR2_596(g25610,g24923,g18127);
  OR2 OR2_597(g31257,g29531,g28253);
  OR2 OR2_598(g25705,g25069,g18744);
  OR2 OR2_599(g28605,g27341,g26302);
  OR2 OR2_600(g33257,g32108,g29519);
  OR2 OR2_601(g32123,g30915,g30919);
  OR2 OR2_602(g33979,g33942,g18361);
  OR2 OR2_603(g33055,g31986,g21976);
  OR2 OR2_604(g16187,g8822,g13486);
  OR2 OR2_605(g25679,g24728,g21836);
  OR2 OR2_606(g33070,g32010,g22114);
  OR2 OR2_607(g33978,g33892,g18356);
  OR2 OR2_608(g25678,g24709,g21835);
  OR2 OR2_609(g26915,g25900,g18230);
  OR2 OR2_610(g33590,g33358,g18470);
  OR2 OR2_611(g15965,g13035,g10675);
  OR2 OR2_612(g28371,g27177,g15847);
  OR4 OR4_18(I30745,g31777,g32321,g32069,g32084);
  OR2 OR2_613(g32230,g30589,g29345);
  OR2 OR2_614(g33986,g33639,g18387);
  OR2 OR2_615(g24252,g22518,g18299);
  OR2 OR2_616(g25686,g24712,g21881);
  OR2 OR2_617(g33384,g32248,g29943);
  OR2 OR2_618(g33067,g31989,g22111);
  OR2 OR2_619(g12768,g7785,g7202);
  OR2 OR2_620(g29250,g28695,g18460);
  OR2 OR2_621(g32992,g32242,g18351);
  OR2 OR2_622(g32391,g31502,g29982);
  OR2 OR2_623(g30455,g30041,g21864);
  OR2 OR2_624(g34455,g34284,g18668);
  OR3 OR3_18(g11372,g490,g482,g8038);
  OR2 OR2_625(g31877,g31278,g21732);
  OR2 OR2_626(g30470,g30165,g21941);
  OR2 OR2_627(g34617,g34526,g18579);
  OR2 OR2_628(g22648,g18987,g15652);
  OR3 OR3_19(I12611,g1500,g1582,g1333);
  OR2 OR2_629(g29296,g28586,g18781);
  OR2 OR2_630(g33019,g32339,g18536);
  OR2 OR2_631(g30201,g23412,g28557);
  OR2 OR2_632(g33018,g32312,g18525);
  OR4 OR4_19(I30761,g32071,g32167,g32067,g32082);
  OR2 OR2_633(g30467,g30185,g21938);
  OR2 OR2_634(g30494,g30209,g21990);
  OR2 OR2_635(g34467,g34341,g18717);
  OR2 OR2_636(g34494,g26849,g34413);
  OR2 OR2_637(g29197,g27187,g27163);
  OR2 OR2_638(g34623,g34525,g18585);
  OR2 OR2_639(g34037,g33803,g18734);
  OR4 OR4_20(I30400,g31021,g30937,g31327,g30614);
  OR2 OR2_640(g27248,g24880,g25953);
  OR2 OR2_641(g30984,g29765,g29755);
  OR2 OR2_642(g27552,g26092,g24676);
  OR2 OR2_643(g31917,g31478,g22003);
  OR2 OR2_644(g30419,g29759,g21803);
  OR2 OR2_645(g31866,g31252,g18142);
  OR2 OR2_646(g30352,g30094,g18340);
  OR2 OR2_647(g27779,g17317,g26694);
  OR2 OR2_648(g25617,g25466,g18189);
  OR2 OR2_649(g24213,g23220,g18186);
  OR3 OR3_20(g23184,g20198,g20185,I22280);
  OR2 OR2_650(g28724,g27491,g16707);
  OR2 OR2_651(g34352,g26079,g34109);
  OR2 OR2_652(g28359,g27151,g15838);
  OR2 OR2_653(g30418,g29751,g21802);
  OR2 OR2_654(g32275,g31210,g29732);
  OR2 OR2_655(g31001,g29360,g28151);
  OR2 OR2_656(g28358,g27149,g15837);
  OR2 OR2_657(g34266,g34076,g18719);
  OR2 OR2_658(g33001,g32282,g18404);
  OR2 OR2_659(g34170,g33790,g19855);
  OR2 OR2_660(g24205,g23006,g18109);
  OR2 OR2_661(g33706,g32412,g33440);
  OR2 OR2_662(g33597,g33344,g18495);
  OR2 OR2_663(g32237,g31153,g29667);
  OR2 OR2_664(g31256,g25983,g29537);
  OR2 OR2_665(g33256,g32107,g29517);
  OR2 OR2_666(g25595,g24835,g21717);
  OR2 OR2_667(g31923,g31763,g22048);
  OR2 OR2_668(g32983,g31990,g18222);
  OR2 OR2_669(g19879,g15841,g13265);
  OR2 OR2_670(g28344,g27136,g15820);
  OR2 OR2_671(g22832,g19354,g15722);
  OR2 OR2_672(g33280,g32141,g29574);
  OR2 OR2_673(g25623,g24552,g18219);
  OR2 OR2_674(g20051,g15936,g13306);
  OR2 OR2_675(g25037,g23103,g19911);
  OR2 OR2_676(g33624,g33371,g18808);
  OR2 OR2_677(g34167,g33786,g19768);
  OR2 OR2_678(g34194,g33811,g33815);
  OR4 OR4_21(g26616,g24881,g24855,g24843,g24822);
  OR2 OR2_679(g19337,g17770,g17785);
  OR2 OR2_680(g28682,g27430,g16635);
  OR2 OR2_681(g29257,g28228,g18600);
  OR4 OR4_22(I23755,g22904,g22927,g22980,g23444);
  OR2 OR2_682(g30524,g30255,g22070);
  OR2 OR2_683(g27233,g25876,g24451);
  OR2 OR2_684(g16800,g13436,g11027);
  OR2 OR2_685(g29496,g28567,g27615);
  OR2 OR2_686(g27182,g25818,g24410);
  OR2 OR2_687(g30401,g29782,g21760);
  OR2 OR2_688(g30477,g30239,g21948);
  OR2 OR2_689(g26305,g24556,g24564);
  OR2 OR2_690(g24350,g23755,g18806);
  OR2 OR2_691(g26809,g24930,g24939);
  OR2 OR2_692(g33066,g32341,g22096);
  OR2 OR2_693(g26900,g26819,g24217);
  OR2 OR2_694(g33231,g32032,g32036);
  OR2 OR2_695(g29741,g28205,g15883);
  OR2 OR2_696(g32130,g30921,g30925);
  OR2 OR2_697(g34022,g33873,g18538);
  OR2 OR2_698(g28134,g27958,g27962);
  OR2 OR2_699(g31876,g31125,g21731);
  OR2 OR2_700(g31885,g31017,g21779);
  OR2 OR2_701(g32362,g29870,g31301);
  OR2 OR2_702(g34616,g34519,g18577);
  OR2 OR2_703(g25589,g21690,g24159);
  OR2 OR2_704(g29801,g25987,g28251);
  OR2 OR2_705(g29735,g28202,g10898);
  OR2 OR2_706(g25588,g21686,g24158);
  OR2 OR2_707(g34305,g25775,g34050);
  OR2 OR2_708(g25836,g25368,g23856);
  OR2 OR2_709(g27026,g26828,g17726);
  OR2 OR2_710(g34254,g34116,g24301);
  OR2 OR2_711(g30466,g30174,g21937);
  OR2 OR2_712(g34809,g33677,g34738);
  OR2 OR2_713(g34900,g34860,g21686);
  OR2 OR2_714(g26733,g10776,g24447);
  OR2 OR2_715(g34466,g34337,g18716);
  OR2 OR2_716(g34808,g34765,g18599);
  OR2 OR2_717(g32222,g31141,g29636);
  OR3 OR3_21(g23771,g21432,g21416,I22912);
  OR2 OR2_718(g26874,I25612,I25613);
  OR2 OR2_719(g34036,g33722,g18715);
  OR2 OR2_720(g30560,g30278,g22131);
  OR2 OR2_721(g34101,g33693,g33700);
  OR2 OR2_722(g31916,g31756,g22002);
  OR2 OR2_723(g34642,g34482,g18725);
  OR2 OR2_724(g25749,g25094,g18800);
  OR2 OR2_725(g25616,g25096,g18172);
  OR2 OR2_726(g28649,g27390,g16597);
  OR2 OR2_727(g33550,g33342,g18338);
  OR2 OR2_728(g32347,g29839,g31273);
  OR2 OR2_729(g33314,g29663,g32174);
  OR2 OR2_730(g31287,g29578,g28292);
  OR2 OR2_731(g15800,g10821,g13242);
  OR2 OR2_732(g32253,g24771,g31207);
  OR2 OR2_733(g25748,g25078,g18799);
  OR2 OR2_734(g33287,g32146,g29586);
  OR2 OR2_735(g34064,g33919,g33922);
  OR2 OR2_736(g30733,g13807,g29773);
  OR2 OR2_737(g31307,g29596,g28311);
  OR2 OR2_738(g33076,g32336,g32446);
  OR2 OR2_739(g34733,g34678,g18651);
  OR2 OR2_740(g26892,g26719,g24198);
  OR2 OR2_741(g25704,g25173,g21925);
  OR2 OR2_742(g22447,g21464,g12761);
  OR2 OR2_743(g33596,g33341,g18494);
  OR2 OR2_744(g33054,g31975,g21975);
  OR2 OR2_745(g32236,g31152,g29664);
  OR2 OR2_746(g8790,I12782,I12783);
  OR2 OR2_747(g32351,g29851,g31281);
  OR2 OR2_748(g32372,g29884,g31314);
  OR2 OR2_749(g34630,g34560,g15117);
  OR2 OR2_750(g34693,g34513,g34310);
  OR2 OR2_751(g24282,g23407,g18657);
  OR2 OR2_752(g26914,g25949,g18227);
  OR2 OR2_753(g29706,g28198,g27208);
  OR2 OR2_754(g8461,g301,g534);
  OR2 OR2_755(g31269,g26024,g29569);
  OR2 OR2_756(g34166,g33785,g19752);
  OR2 OR2_757(g34009,g33863,g18477);
  OR2 OR2_758(g19336,g17769,g14831);
  OR2 OR2_759(g26907,g26513,g24224);
  OR2 OR2_760(g29256,g28597,g18533);
  OR2 OR2_761(g31773,g30044,g30056);
  OR4 OR4_23(I30399,g29385,g31376,g30735,g30825);
  OR2 OR2_762(g31268,g29552,g28266);
  OR2 OR2_763(g32264,g31187,g29711);
  OR2 OR2_764(g34008,g33849,g18476);
  OR2 OR2_765(g29280,g28530,g18742);
  OR2 OR2_766(g33268,g32116,g29538);
  OR2 OR2_767(g30476,g30229,g21947);
  OR2 OR2_768(g30485,g30166,g21981);
  OR2 OR2_769(g29300,g28666,g18796);
  OR2 OR2_770(g31670,g29937,g28573);
  OR2 OR2_771(g8904,g1779,g1798);
  OR4 OR4_24(I31863,g33506,g33507,g33508,g33509);
  OR2 OR2_772(g30555,g30227,g22126);
  OR2 OR2_773(g30454,g29909,g21863);
  OR2 OR2_774(g34454,g34414,g18667);
  OR2 OR2_775(g25733,g25108,g18778);
  OR3 OR3_22(g13091,g329,g319,g10796);
  OR2 OR2_776(g22591,g18893,g18909);
  OR2 OR2_777(g27133,g25788,g24392);
  OR2 OR2_778(g28719,g27485,g16703);
  OR4 OR4_25(g28191,g27217,g27210,g27186,g27162);
  OR2 OR2_779(g31930,g31769,g22094);
  OR2 OR2_780(g32209,g31122,g29599);
  OR2 OR2_781(g33993,g33646,g18413);
  OR2 OR2_782(g25630,g24532,g18263);
  OR2 OR2_783(g28718,g27483,g16702);
  OR2 OR2_784(g25693,g24627,g18707);
  OR2 OR2_785(g29231,g28301,g18229);
  OR2 OR2_786(g33694,g32402,g33429);
  OR2 OR2_787(g32208,g31120,g29584);
  OR2 OR2_788(g33965,g33805,g18179);
  OR4 OR4_26(I12783,g4204,g4207,g4210,g4180);
  OR2 OR2_789(g25665,g24708,g21790);
  OR2 OR2_790(g34239,g32845,g33957);
  OR2 OR2_791(g34238,g32780,g33956);
  OR2 OR2_792(g23345,g19735,g16203);
  OR2 OR2_793(g26883,g26670,g24189);
  OR4 OR4_27(I23162,g19919,g19968,g20014,g20841);
  OR2 OR2_794(g33619,g33359,g18758);
  OR2 OR2_795(g33557,g33331,g18363);
  OR2 OR2_796(g29763,g28217,g22762);
  OR2 OR2_797(g30382,g30137,g18498);
  OR2 OR2_798(g30519,g30264,g22040);
  OR2 OR2_799(g33618,g33353,g18757);
  OR2 OR2_800(g28389,g27206,g15860);
  OR2 OR2_801(g30176,g23392,g28531);
  OR2 OR2_802(g28045,g27378,g18141);
  OR2 OR2_803(g30092,g28466,g16699);
  OR2 OR2_804(g31279,g29571,g29579);
  OR2 OR2_805(g24249,g22624,g18294);
  OR2 OR2_806(g33279,g32140,g29573);
  OR2 OR2_807(g25712,g25126,g21963);
  OR2 OR2_808(g28099,g27992,g22043);
  OR2 OR2_809(g30518,g30254,g22039);
  OR3 OR3_23(I22280,g20271,g20150,g20134);
  OR2 OR2_810(g28388,g27204,g15859);
  OR2 OR2_811(g16430,g182,g13657);
  OR2 OR2_812(g28701,g27455,g16669);
  OR2 OR2_813(g24248,g22710,g18286);
  OR2 OR2_814(g33278,g32139,g29572);
  OR2 OR2_815(g12925,g8928,g10511);
  OR2 OR2_816(g28777,g27539,g16807);
  OR2 OR2_817(g28534,g27292,g26204);
  OR2 OR2_818(g28098,g27683,g22016);
  OR2 OR2_819(g32346,g29838,g31272);
  OR2 OR2_820(g34637,g34478,g18694);
  OR2 OR2_821(g24204,g22990,g18108);
  OR2 OR2_822(g33286,g32145,g29585);
  OR2 OR2_823(g31468,g29641,g29656);
  OR2 OR2_824(g31306,g29595,g29610);
  OR4 OR4_28(I31873,g33524,g33525,g33526,g33527);
  OR2 OR2_825(g33039,g32187,g24312);
  OR2 OR2_826(g29480,g28115,g22172);
  OR2 OR2_827(g27742,g17292,g26673);
  OR2 OR2_828(g22318,g21394,g17783);
  OR2 OR2_829(g25594,g24772,g21708);
  OR2 OR2_830(g33038,g32184,g24311);
  OR2 OR2_831(g29287,g28555,g18760);
  OR2 OR2_832(g29307,g28706,g18814);
  OR2 OR2_833(g28140,I26643,I26644);
  OR2 OR2_834(g26349,g24630,g13409);
  OR2 OR2_835(g33601,g33422,g18508);
  OR2 OR2_836(g25941,g24416,g22219);
  OR3 OR3_24(g33187,g32014,I30740,I30741);
  OR2 OR2_837(g33975,g33860,g18346);
  OR2 OR2_838(g27429,g25969,g24589);
  OR2 OR2_839(g26906,g26423,g24223);
  OR2 OR2_840(g25675,g24769,g21832);
  OR2 OR2_841(g29243,g28657,g18358);
  OR2 OR2_842(g26348,g8466,g24609);
  OR2 OR2_843(g30501,g29327,g22018);
  OR2 OR2_844(g28061,g27287,g21735);
  OR2 OR2_845(g34729,g34666,g18270);
  OR2 OR2_846(g32408,g31541,g30073);
  OR2 OR2_847(g30439,g29761,g21848);
  OR2 OR2_848(g34728,g34661,g18214);
  OR2 OR2_849(g34439,g34344,g18181);
  OR2 OR2_850(g29269,g28249,g18634);
  OR2 OR2_851(g25637,g24618,g18307);
  OR2 OR2_852(g24233,g22590,g18236);
  OR2 OR2_853(g25935,g24402,g22208);
  OR2 OR2_854(g30438,g29890,g21847);
  OR2 OR2_855(g19525,g7696,g16811);
  OR2 OR2_856(g19488,g16965,g14148);
  OR2 OR2_857(g34438,g34348,g18150);
  OR2 OR2_858(g29268,g28343,g18625);
  OR4 OR4_29(I25613,g25571,g25572,g25573,g25574);
  OR2 OR2_859(g31884,g31290,g21778);
  OR2 OR2_860(g33791,g33379,g32430);
  OR2 OR2_861(g30349,g30051,g18333);
  OR2 OR2_862(g34349,g26019,g34104);
  OR3 OR3_25(g8417,g1056,g1116,I12583);
  OR2 OR2_863(g30348,g30083,g18329);
  OR2 OR2_864(g22645,g18982,g15633);
  OR2 OR2_865(g34906,g34857,g21694);
  OR2 OR2_866(g29734,g28201,g15872);
  OR2 OR2_867(g30304,g28255,g27259);
  OR2 OR2_868(g33015,g32343,g18507);
  OR2 OR2_869(g34622,g34520,g18584);
  OR2 OR2_870(g25729,g25091,g22012);
  OR4 OR4_30(g26636,g24897,g24884,g24858,g24846);
  OR2 OR2_871(g28629,g27371,g16532);
  OR2 OR2_872(g25577,g24143,g24144);
  OR3 OR3_26(g28220,g23495,I26741,I26742);
  OR2 OR2_873(g25728,g25076,g22011);
  OR2 OR2_874(g28628,g27370,g16531);
  OR2 OR2_875(g33556,g33329,g18362);
  OR2 OR2_876(g24212,g23280,g18155);
  OR2 OR2_877(g26963,g26306,g24308);
  OR2 OR2_878(g33580,g33330,g18442);
  OR2 OR2_879(g29487,g25815,g28133);
  OR2 OR2_880(g23795,g20203,g16884);
  OR2 OR2_881(g28071,g27085,g21873);
  OR2 OR2_882(g29502,g28139,g25871);
  OR2 OR2_883(g27533,g26078,g24659);
  OR4 OR4_31(I29351,g29328,g29323,g29316,g30316);
  OR2 OR2_884(g28591,g27332,g26286);
  OR2 OR2_885(g25906,g25559,g24014);
  OR2 OR2_886(g28776,g27538,g13974);
  OR2 OR2_887(g30415,g29843,g21799);
  OR2 OR2_888(g30333,g29834,g21699);
  OR2 OR2_889(g34636,g34476,g18693);
  OR2 OR2_890(g22547,g16855,g20215);
  OR2 OR2_891(g29279,g28442,g18741);
  OR2 OR2_892(g31922,g31525,g22047);
  OR2 OR2_893(g32982,g31948,g18208);
  OR2 OR2_894(g33321,g29712,g32182);
  OR2 OR2_895(g25622,g24546,g18217);
  OR2 OR2_896(g29278,g28626,g18740);
  OR2 OR2_897(g19267,g17752,g17768);
  OR2 OR2_898(g22226,g21333,g17655);
  OR2 OR2_899(g24433,g10878,g22400);
  OR2 OR2_900(g20148,g16128,g13393);
  OR2 OR2_901(g29286,g28542,g18759);
  OR2 OR2_902(g27232,g25874,g24450);
  OR2 OR2_903(g7404,g933,g939);
  OR2 OR2_904(g29306,g28689,g18813);
  OR4 OR4_32(g28172,g27469,g27440,g27416,g27395);
  OR2 OR2_905(g33685,g32396,g33423);
  OR2 OR2_906(g7764,g2999,g2932);
  OR3 OR3_27(g33953,g33487,I31848,I31849);
  OR2 OR2_907(g24343,g23724,g18773);
  OR2 OR2_908(g26921,g25955,g18285);
  OR2 OR2_909(g25653,g24664,g18602);
  OR2 OR2_910(g32390,g31501,g29979);
  OR2 OR2_911(g27261,g24544,g25996);
  OR2 OR2_912(g30484,g30154,g21980);
  OR2 OR2_913(g30554,g30216,g22125);
  OR2 OR2_914(g22490,g21513,g12795);
  OR3 OR3_28(g13820,g11184,g9187,g12527);
  OR2 OR2_915(g26813,g24940,g24949);
  OR4 OR4_33(g15727,g13383,g13345,g13333,g11010);
  OR2 OR2_916(g25636,g24507,g18305);
  OR2 OR2_917(g30609,g13633,g29742);
  OR2 OR2_918(g34609,g34503,g18563);
  OR2 OR2_919(g28420,g27222,g13290);
  OR2 OR2_920(g30608,g13604,g29736);
  OR2 OR2_921(g28319,g27115,g15807);
  OR2 OR2_922(g30115,g28489,g11449);
  OR2 OR2_923(g29143,g27650,g17146);
  OR2 OR2_924(g34608,g34568,g15082);
  OR4 OR4_34(g17490,g14364,g14337,g11958,I18421);
  OR2 OR2_925(g26805,g10776,g24478);
  OR2 OR2_926(g31762,g30011,g30030);
  OR2 OR2_927(g23358,g19746,g16212);
  OR4 OR4_35(I30760,g31778,g32295,g32046,g32050);
  OR2 OR2_928(g31964,g31654,g14544);
  OR2 OR2_929(g33964,g33817,g18146);
  OR2 OR2_930(g25664,g24681,g21789);
  OR2 OR2_931(g28059,g27042,g18276);
  OR2 OR2_932(g29791,g28233,g22859);
  OR2 OR2_933(g16021,g13047,g10706);
  OR2 OR2_934(g26934,g26845,g18556);
  OR2 OR2_935(g28058,g27235,g18268);
  OR2 OR2_936(g29168,g27658,g26613);
  OR2 OR2_937(g33587,g33363,g18463);
  OR2 OR2_938(g24896,g22863,g19684);
  OR2 OR2_939(g34799,g34751,g18578);
  OR2 OR2_940(g25585,g21674,g24155);
  OR2 OR2_941(g25576,g24141,g24142);
  OR2 OR2_942(g29479,g28113,g28116);
  OR2 OR2_943(g34798,g34754,g18575);
  OR2 OR2_944(g31909,g31750,g21956);
  OR2 OR2_945(g28044,g27256,g18130);
  OR2 OR2_946(g33543,g33106,g18281);
  OR2 OR2_947(g19595,g17149,g14218);
  OR2 OR2_948(g29478,g28111,g22160);
  OR2 OR2_949(g19467,g16896,g14097);
  OR2 OR2_950(g25609,g24915,g18126);
  OR2 OR2_951(g34805,g34748,g18594);
  OR2 OR2_952(g31908,g31519,g21955);
  OR2 OR2_953(g33000,g32270,g18403);
  OR2 OR2_954(g29486,g28537,g27595);
  OR2 OR2_955(g32252,g31183,g31206);
  OR2 OR2_956(g25608,g24643,g18120);
  OR2 OR2_957(g33569,g33415,g18402);
  OR2 OR2_958(g30732,g13778,g29762);
  OR2 OR2_959(g27271,g24547,g26053);
  OR3 OR3_29(I18495,g14539,g14515,g14449);
  OR2 OR2_960(g34732,g34686,g18593);
  OR2 OR2_961(g26329,g8526,g24609);
  OR2 OR2_962(g33568,g33409,g18395);
  OR2 OR2_963(g25745,g25150,g22060);
  OR2 OR2_964(g29223,g28341,g18131);
  OR2 OR2_965(g26328,g1183,g24591);
  OR2 OR2_966(g28562,g27313,g26251);
  OR2 OR2_967(g14844,g10776,g8703);
  OR2 OR2_968(g34761,g34679,g34506);
  OR2 OR2_969(g28699,g27452,g16667);
  OR4 OR4_36(g27031,g26213,g26190,g26166,g26148);
  OR2 OR2_970(g33123,g31962,g30577);
  OR4 OR4_37(I30755,g30564,g32303,g32049,g32055);
  OR2 OR2_971(g28698,g27451,g16666);
  OR2 OR2_972(g31751,g29975,g29990);
  OR2 OR2_973(g31772,g30035,g28654);
  OR2 OR2_974(g30400,g29766,g21759);
  OR2 OR2_975(g33974,g33846,g18345);
  OR2 OR2_976(g30214,g23424,g28572);
  OR2 OR2_977(g34013,g33901,g18488);
  OR4 OR4_38(g25805,g25453,g25414,g25374,g25331);
  OR2 OR2_978(g25674,g24755,g21831);
  OR2 OR2_979(g31293,g29582,g28299);
  OR2 OR2_980(g33293,g32151,g29602);
  OR2 OR2_981(g30539,g30267,g22085);
  OR2 OR2_982(g34207,g33835,g33304);
  OR2 OR2_983(g22659,g19062,g15673);
  OR2 OR2_984(g22625,g18910,g18933);
  OR2 OR2_985(g25732,g25201,g22017);
  OR2 OR2_986(g34005,g33883,g18454);
  OR2 OR2_987(g28632,g27373,g16535);
  OR2 OR2_988(g33265,g32113,g29530);
  OR2 OR2_989(g30538,g30256,g22084);
  OR2 OR2_990(g29373,g13832,g28453);
  OR4 OR4_39(I30262,g31672,g31710,g31021,g30937);
  OR2 OR2_991(g33992,g33900,g18408);
  OR2 OR2_992(g25761,g25152,g18812);
  OR2 OR2_993(g28661,g27406,g16611);
  OR2 OR2_994(g28403,g27214,g13282);
  OR2 OR2_995(g22644,g18981,g15632);
  OR4 OR4_40(I12782,g4188,g4194,g4197,g4200);
  OR2 OR2_996(g33579,g33357,g18437);
  OR2 OR2_997(g14044,g10776,g8703);
  OR2 OR2_998(g28715,g27480,g16700);
  OR4 OR4_41(I30718,g32348,g32356,g32097,g32020);
  OR2 OR2_999(g33578,g33410,g18433);
  OR2 OR2_1000(g31014,g29367,g28160);
  OR2 OR2_1001(g27225,g2975,g26364);
  OR2 OR2_1002(g33014,g32305,g18499);
  OR2 OR2_1003(g23770,g20188,g16868);
  OR2 OR2_1004(g26882,g26650,g24188);
  OR2 OR2_1005(g28551,g27305,g26234);
  OR2 OR2_1006(g31007,g29364,g28159);
  OR2 OR2_1007(g27258,g25905,g15749);
  OR2 OR2_1008(g34100,g33690,g33697);
  OR2 OR2_1009(g33586,g33416,g18459);
  OR2 OR2_1010(g33007,g32331,g18455);
  OR2 OR2_1011(g25539,g23531,g20628);
  OR2 OR2_1012(g13662,g10896,g10917);
  OR2 OR2_1013(g34235,g32585,g33953);
  OR2 OR2_1014(g27244,g24652,g25995);
  OR2 OR2_1015(g28490,g27262,g16185);
  OR2 OR2_1016(g33116,g32403,g32411);
  OR2 OR2_1017(g33615,g33113,g21871);
  OR2 OR2_1018(g23262,g19661,g16126);
  OR2 OR2_1019(g21899,g20162,g15113);
  OR2 OR2_1020(g30515,g30223,g22036);
  OR2 OR2_1021(g30414,g30002,g21794);
  OR2 OR2_1022(g28385,g27201,g15857);
  OR2 OR2_1023(g33041,g32189,g24323);
  OR2 OR2_1024(g28297,g27096,g15785);
  OR2 OR2_1025(g21898,g20152,g15112);
  OR2 OR2_1026(g34882,g34876,g18659);
  OR2 OR2_1027(g28103,g27696,g22097);
  OR2 OR2_1028(g24245,g22849,g18256);
  OR2 OR2_1029(g33275,g32127,g29564);
  OR2 OR2_1030(g28095,g27674,g21970);
  OR2 OR2_1031(g30407,g29794,g21766);
  OR2 OR2_1032(g34407,g34185,g25124);
  OR2 OR2_1033(g27970,g26514,g25050);
  OR2 OR2_1034(g31465,g26156,g29647);
  OR2 OR2_1035(g26759,g24468,g7511);
  OR2 OR2_1036(g26725,g24457,g10719);
  OR2 OR2_1037(g28671,g27413,g16619);
  OR2 OR2_1038(g33983,g33877,g18373);
  OR2 OR2_1039(g22707,g20559,g17156);
  OR2 OR2_1040(g33035,g32019,g21872);
  OR2 OR2_1041(g27886,g14438,g26759);
  OR2 OR2_1042(g25683,g24669,g18641);
  OR2 OR2_1043(g29242,g28674,g18354);
  OR2 OR2_1044(g26082,g2898,g24561);
  OR2 OR2_1045(g11380,g8583,g8530);
  OR2 OR2_1046(g30441,g29787,g21850);
  OR2 OR2_1047(g34441,g34381,g18540);
  OR2 OR2_1048(g24232,g22686,g18228);
  OR2 OR2_1049(g34206,g33834,g33836);
  OR2 OR2_1050(g26940,g25908,g21886);
  OR4 OR4_42(I25612,g25567,g25568,g25569,g25570);
  OR2 OR2_1051(g34725,g34700,g18183);
  OR2 OR2_1052(g24261,g22862,g18314);
  OR2 OR2_1053(g29230,g28107,g18202);
  OR2 OR2_1054(g27458,g24590,g25989);
  OR2 OR2_1055(g29293,g28570,g18777);
  OR2 OR2_1056(g30114,g28488,g16761);
  OR2 OR2_1057(g30435,g30025,g21840);
  OR2 OR2_1058(g29265,g28318,g18620);
  OR2 OR2_1059(g28546,g27302,g26231);
  OR2 OR2_1060(g28089,g27269,g18731);
  OR2 OR2_1061(g23251,g19637,g16098);
  OR2 OR2_1062(g28211,g27029,g27034);
  OR2 OR2_1063(g34107,g33710,g33121);
  OR2 OR2_1064(g19555,g15672,g13030);
  OR2 OR2_1065(g28088,g27264,g18729);
  OR2 OR2_1066(g30345,g29644,g18302);
  OR2 OR2_1067(g30399,g29757,g21758);
  OR2 OR2_1068(g34849,g34842,g18154);
  OR2 OR2_1069(g34399,g34178,g25067);
  OR2 OR2_1070(g25584,g21670,g24154);
  OR2 OR2_1071(g28497,g27267,g16199);
  OR2 OR2_1072(g33006,g32291,g18447);
  OR2 OR2_1073(g30398,g29749,g21757);
  OR2 OR2_1074(g26962,g26295,g24307);
  OR2 OR2_1075(g26361,g24674,g22991);
  OR2 OR2_1076(g23997,g20602,g17191);
  OR2 OR2_1077(g30141,g28499,g16844);
  OR2 OR2_1078(g34804,g34740,g18591);
  OR2 OR2_1079(g28700,g27454,g16668);
  OR2 OR2_1080(g25759,g25166,g22106);
  OR2 OR2_1081(g28659,g27404,g16610);
  OR2 OR2_1082(g25725,g25127,g22008);
  OR2 OR2_1083(g28625,g27363,g26324);
  OR2 OR2_1084(g14888,g10776,g8703);
  OR2 OR2_1085(g32357,g29865,g31296);
  OR2 OR2_1086(g27159,g25814,g12953);
  OR2 OR2_1087(g27532,g16176,g26084);
  OR2 OR2_1088(g25758,g25151,g22105);
  OR2 OR2_1089(g34263,g34078,g18699);
  OR2 OR2_1090(g34332,g34071,g33723);
  OR2 OR2_1091(g33703,g32410,g33434);
  OR2 OR2_1092(g28296,g27095,g15784);
  OR2 OR2_1093(g31253,g25980,g29533);
  OR2 OR2_1094(g27561,g26100,g24702);
  OR2 OR2_1095(g33253,g32103,g29511);
  OR2 OR2_1096(g25744,g25129,g22059);
  OR2 OR2_1097(g28644,g27387,g16593);
  OR2 OR2_1098(g30406,g29783,g21765);
  OR2 OR2_1099(g24432,g23900,g21361);
  OR2 OR2_1100(g30361,g30109,g18391);
  OR2 OR2_1101(g34406,g34184,g25123);
  OR2 OR2_1102(g24271,g23451,g18628);
  OR2 OR2_1103(g33600,g33418,g18501);
  OR2 OR2_1104(g25940,g24415,g22218);
  OR2 OR2_1105(g31781,g30058,g30069);
  OR3 OR3_30(g23162,g20184,g20170,I22267);
  OR2 OR2_1106(g33236,g32044,g32045);
  OR2 OR2_1107(g30500,g29326,g21996);
  OR2 OR2_1108(g29275,g28165,g21868);
  OR2 OR2_1109(g28060,g27616,g18532);
  OR3 OR3_31(g33952,g33478,I31843,I31844);
  OR2 OR2_1110(g24342,g23691,g18772);
  OR2 OR2_1111(g25652,g24777,g21747);
  OR2 OR2_1112(g26947,g26394,g24285);
  OR2 OR2_1113(g8905,g2204,g2223);
  OR2 OR2_1114(g29237,g28185,g18289);
  OR2 OR2_1115(g28527,g27286,g26182);
  OR2 OR2_1116(g33063,g31988,g22066);
  OR2 OR2_1117(g34004,g33879,g18453);
  OR2 OR2_1118(g26951,g26390,g24289);
  OR2 OR2_1119(g26972,g26780,g25229);
  OR2 OR2_1120(g31873,g31270,g21728);
  OR2 OR2_1121(g19501,g16986,g14168);
  OR2 OR2_1122(g34613,g34515,g18567);
  OR2 OR2_1123(g32249,g31169,g29687);
  OR2 OR2_1124(g30605,g29529,g29520);
  OR2 OR2_1125(g27289,g25925,g25927);
  OR2 OR2_1126(g34273,g27765,g34203);
  OR2 OR2_1127(g34605,g34566,g15077);
  OR2 OR2_1128(g18879,g17365,g14423);
  OR2 OR2_1129(g28581,g27329,g26276);
  OR2 OR2_1130(g27224,g25870,g15678);
  OR2 OR2_1131(g30463,g30140,g21934);
  OR2 OR2_1132(g27571,g26127,g24723);
  OR2 OR2_1133(g28707,g27461,g16673);
  OR2 OR2_1134(g34463,g34338,g18686);
  OR2 OR2_1135(g23825,g20705,g20781);
  OR2 OR2_1136(g30371,g30099,g18445);
  OR2 OR2_1137(g28818,g27549,g13998);
  OR2 OR2_1138(g34033,g33821,g18708);
  OR2 OR2_1139(g34234,g32520,g33952);
  OR2 OR2_1140(g28055,g27560,g18190);
  OR2 OR2_1141(g33542,g33102,g18265);
  OR2 OR2_1142(g33021,g32302,g21749);
  OR2 OR2_1143(g24259,g23008,g18312);
  OR2 OR2_1144(g28070,g27050,g21867);
  OR2 OR2_1145(g31913,g31485,g21999);
  OR2 OR2_1146(g18994,g16303,g13632);
  OR2 OR2_1147(g24471,g10999,g22450);
  OR2 OR2_1148(g34795,g34753,g18572);
  OR2 OR2_1149(g25613,g25181,g18140);
  OR2 OR2_1150(g24258,g22851,g18311);
  OR2 OR2_1151(g33614,g33249,g18650);
  OR4 OR4_43(g17511,g14396,g14365,g11976,I18452);
  OR2 OR2_1152(g32999,g32337,g18401);
  OR2 OR2_1153(g33607,g33091,g18526);
  OR2 OR2_1154(g31905,g31746,g21952);
  OR2 OR2_1155(g31320,g26125,g29632);
  OR2 OR2_1156(g30514,g30211,g22035);
  OR2 OR2_1157(g32380,g29907,g31467);
  OR2 OR2_1158(g31274,g29565,g28280);
  OR2 OR2_1159(g25605,g24743,g18116);
  OR2 OR2_1160(g29222,g28252,g18105);
  OR2 OR2_1161(g24244,g23349,g18255);
  OR2 OR2_1162(g33274,g32126,g29563);
  OR2 OR2_1163(g30507,g30190,g22028);
  OR2 OR2_1164(g32998,g32300,g18393);
  OR2 OR2_1165(g28094,g27673,g21959);
  OR2 OR2_1166(g28067,g27309,g21827);
  OR2 OR2_1167(g33593,g33417,g18482);
  OR2 OR2_1168(g26789,g10776,g24471);
  OR2 OR2_1169(g32233,g31150,g29661);
  OR2 OR2_1170(g12954,g12186,g9906);
  OR2 OR2_1171(g23319,g19717,g16193);
  OR2 OR2_1172(g30421,g29784,g21805);
  OR2 OR2_1173(g33565,g33338,g18389);
  OR2 OR2_1174(g34421,g27686,g34198);
  OR2 OR2_1175(g26359,g24651,g22939);
  OR2 OR2_1176(g28735,g27510,g16737);
  OR2 OR2_1177(g23318,g19716,g16192);
  OR2 OR2_1178(g30163,g23381,g28523);
  OR2 OR2_1179(g33034,g32340,g21844);
  OR2 OR2_1180(g26920,g25865,g18283);
  OR2 OR2_1181(g34012,g33886,g18480);
  OR2 OR2_1182(g29253,g28697,g18490);
  OR2 OR2_1183(g24879,g21465,g24009);
  OR2 OR2_1184(g33292,g32150,g29601);
  OR2 OR2_1185(g26946,g26389,g24284);
  OR2 OR2_1186(g30541,g30281,g22087);
  OR2 OR2_1187(g30473,g30196,g21944);
  OR2 OR2_1188(g24337,g23540,g18754);
  OR2 OR2_1189(g27489,g24608,g26022);
  OR2 OR2_1190(g29236,g28313,g18287);
  OR2 OR2_1191(g28526,g27285,g26178);
  OR2 OR2_1192(g26344,g2927,g25010);
  OR2 OR2_1193(g27016,g26821,g14585);
  OR2 OR2_1194(g30359,g30075,g18385);
  OR2 OR2_1195(g34724,g34702,g18152);
  OR2 OR2_1196(g28402,g27213,g15873);
  OR2 OR2_1197(g30535,g30225,g22081);
  OR2 OR2_1198(g30434,g30024,g21818);
  OR2 OR2_1199(g19576,g17138,g14202);
  OR2 OR2_1200(g30358,g30108,g18381);
  OR2 OR2_1201(g34535,g34309,g34073);
  OR2 OR2_1202(g29264,g28248,g18618);
  OR2 OR2_1203(g29790,g25975,g28242);
  OR2 OR2_1204(g16928,g13525,g11127);
  OR2 OR2_1205(g27544,g26087,g24671);
  OR3 OR3_32(g33164,g32203,I30727,I30728);
  OR2 OR2_1206(g17268,g9220,g14387);
  OR2 OR2_1207(g24919,g21606,g22143);
  OR2 OR2_1208(g30344,g29630,g18298);
  OR2 OR2_1209(g31891,g31305,g21824);
  OR2 OR2_1210(g28077,g27120,g21879);
  OR2 OR2_1211(g33891,g33264,g33269);
  OR2 OR2_1212(g31474,g29668,g13583);
  OR2 OR2_1213(g33575,g33086,g18420);
  OR2 OR2_1214(g24444,g10890,g22400);
  OR2 OR2_1215(g30291,g28672,g27685);
  OR2 OR2_1216(g25789,g25285,g14543);
  OR2 OR2_1217(g32387,g31489,g29952);
  OR2 OR2_1218(g25724,g25043,g22007);
  OR2 OR2_1219(g28688,g27435,g16639);
  OR2 OR2_1220(g33537,g33244,g21716);
  OR2 OR2_1221(g22487,g21512,g12794);
  OR2 OR2_1222(g28102,g27995,g22089);
  OR2 OR2_1223(g33283,g31995,g30318);
  OR2 OR2_1224(g27383,g24569,g25961);
  OR2 OR2_1225(g33606,g33369,g18522);
  OR2 OR2_1226(g31303,g29592,g29606);
  OR2 OR2_1227(g33303,g32159,g29638);
  OR2 OR2_1228(g34029,g33798,g18703);
  OR2 OR2_1229(g26927,g26711,g18539);
  OR2 OR2_1230(g30506,g30179,g22027);
  OR2 OR2_1231(g28066,g27553,g21819);
  OR2 OR2_1232(g21895,g20135,g15108);
  OR2 OR2_1233(g34028,g33720,g18684);
  OR2 OR2_1234(g32368,g29881,g31310);
  OR2 OR2_1235(g33982,g33865,g18372);
  OR2 OR2_1236(g25682,g24658,g18640);
  OR2 OR2_1237(g29274,g28360,g18642);
  OR2 OR2_1238(g24561,I23755,I23756);
  OR2 OR2_1239(g24353,g23682,g18822);
  OR2 OR2_1240(g26903,g26388,g24220);
  OR2 OR2_1241(g35000,g34953,g34999);
  OR2 OR2_1242(g11737,g8359,g8292);
  OR2 OR2_1243(g9012,g2047,g2066);
  OR2 OR2_1244(g26755,g10776,g24457);
  OR2 OR2_1245(g28511,g27272,g16208);
  OR2 OR2_1246(g32229,g31148,g29652);
  OR2 OR2_1247(g26770,g24471,g10732);
  OR2 OR2_1248(g24336,g24012,g18753);
  OR2 OR2_1249(g27837,g17401,g26725);
  OR2 OR2_1250(g33390,g32276,g29968);
  OR2 OR2_1251(g32228,g31147,g29651);
  OR2 OR2_1252(g25760,g25238,g22109);
  OR2 OR2_1253(g29292,g28556,g18776);
  OR2 OR2_1254(g34649,g33111,g34492);
  OR2 OR2_1255(g34240,g32910,g33958);
  OR2 OR2_1256(g30491,g30178,g21987);
  OR2 OR2_1257(g34903,g34859,g21690);
  OR2 OR2_1258(g23297,g19692,g16178);
  OR2 OR2_1259(g34604,g34563,g15076);
  OR2 OR2_1260(g26899,g26844,g18199);
  OR2 OR2_1261(g30563,g29347,g22134);
  OR2 OR2_1262(g26898,g26387,g18194);
  OR2 OR2_1263(g28085,g27263,g18700);
  OR2 OR2_1264(g28076,g27098,g21878);
  OR2 OR2_1265(g28721,g27488,g16705);
  OR2 OR2_1266(g28596,g27336,g26291);
  OR2 OR2_1267(g28054,g27723,g18170);
  OR2 OR2_1268(g33553,g33403,g18350);
  OR2 OR2_1269(g15803,g12924,g10528);
  OR2 OR2_1270(g22217,g21302,g17617);
  OR2 OR2_1271(g33949,g32446,g33459);
  OR2 OR2_1272(g31326,g29627,g29640);
  OR2 OR2_1273(g32386,g31488,g29949);
  OR2 OR2_1274(g30395,g29841,g21754);
  OR2 OR2_1275(g34794,g34746,g18571);
  OR2 OR2_1276(g25649,g24654,g21742);
  OR4 OR4_44(I26644,g27057,g27044,g27039,g27032);
  OR4 OR4_45(g27037,g26236,g26218,g26195,g26171);
  OR2 OR2_1277(g34262,g34075,g18697);
  OR2 OR2_1278(g33536,g33241,g21715);
  OR2 OR2_1279(g33040,g32164,g24313);
  OR2 OR2_1280(g33948,g32442,g33458);
  OR2 OR2_1281(g25648,g24644,g21741);
  OR2 OR2_1282(g28773,g27535,g16803);
  OR2 OR2_1283(g31757,g29992,g30010);
  OR2 OR2_1284(g31904,g31780,g21923);
  OR2 OR2_1285(g34633,g34481,g18690);
  OR2 OR2_1286(g25604,g24717,g18115);
  OR2 OR2_1287(g25755,g25192,g22102);
  OR2 OR2_1288(g33621,g33365,g18775);
  OR2 OR2_1289(g34719,g34701,g18133);
  OR2 OR2_1290(g28180,g20242,g27511);
  OR2 OR2_1291(g28670,g27412,g16618);
  OR2 OR2_1292(g26926,g26633,g18531);
  OR2 OR2_1293(g32429,g30318,g31794);
  OR2 OR2_1294(g30521,g29331,g22042);
  OR2 OR2_1295(g14511,g10685,g546);
  OR2 OR2_1296(g33564,g33332,g18388);
  OR2 OR2_1297(g26099,g24506,g22538);
  OR2 OR2_1298(g29283,g28627,g18746);
  OR2 OR2_1299(g28734,g27508,g16736);
  OR2 OR2_1300(g28335,g27132,g15818);
  OR2 OR2_1301(g29303,g28703,g18801);
  OR2 OR2_1302(g24374,g19345,g24004);
  OR2 OR2_1303(g30440,g29771,g21849);
  OR2 OR2_1304(g34440,g34364,g24226);
  OR2 OR2_1305(g25767,g25207,g12015);
  OR2 OR2_1306(g28667,g27410,g16616);
  OR2 OR2_1307(g33062,g31977,g22065);
  OR2 OR2_1308(g22531,g20773,g20922);
  OR2 OR2_1309(g27589,g26177,g24763);
  OR2 OR2_1310(g16448,g13287,g10934);
  OR2 OR2_1311(g30389,g29969,g18554);
  OR2 OR2_1312(g24260,g23373,g18313);
  OR2 OR2_1313(g27524,g26050,g24649);
  OR2 OR2_1314(g25633,g24420,g18282);
  OR2 OR2_1315(g31872,g31524,g18535);
  OR2 OR2_1316(g24842,g7804,g22669);
  OR2 OR2_1317(g30388,g30023,g18534);
  OR2 OR2_1318(g34612,g34514,g18566);
  OR2 OR2_1319(g25719,g25089,g18761);
  OR2 OR2_1320(g28619,g27358,g16517);
  OR2 OR2_1321(g34099,g33684,g33689);
  OR2 OR2_1322(g30534,g30213,g22080);
  OR2 OR2_1323(g19441,g15507,g12931);
  OR2 OR2_1324(g25718,g25187,g21971);
  OR2 OR2_1325(g28618,g27357,g16516);
  OR2 OR2_1326(g34251,g34157,g18147);
  OR2 OR2_1327(g28279,g27087,g25909);
  OR2 OR2_1328(g26766,g10776,g24460);
  OR2 OR2_1329(g30462,g30228,g21933);
  OR2 OR2_1330(g23296,g19691,g16177);
  OR2 OR2_1331(g34462,g34334,g18685);
  OR2 OR2_1332(g28286,g27090,g15757);
  OR2 OR2_1333(g32245,g31167,g29684);
  OR2 OR2_1334(g34032,g33816,g18706);
  OR2 OR2_1335(g28306,g27104,g15794);
  OR2 OR2_1336(g33574,g33362,g18416);
  OR2 OR2_1337(g33047,g31944,g21927);
  OR4 OR4_46(I26741,g22881,g22905,g22928,g27402);
  OR2 OR2_1338(g31912,g31752,g21998);
  OR2 OR2_1339(g31311,g26103,g29618);
  OR2 OR2_1340(g23197,g19571,g15966);
  OR2 OR2_1341(g25612,g24941,g18132);
  OR2 OR2_1342(g28815,g27546,g16842);
  OR2 OR2_1343(g29483,g25801,g28130);
  OR2 OR2_1344(g16811,g8690,g13914);
  OR2 OR2_1345(g25701,g25054,g21920);
  OR4 OR4_47(I30055,g31070,g31170,g30614,g30673);
  OR2 OR2_1346(g24705,g2890,g23267);
  OR2 OR2_1347(g33051,g32316,g21958);
  OR2 OR2_1348(g24255,g22835,g18308);
  OR2 OR2_1349(g33592,g33412,g18475);
  OR2 OR2_1350(g30360,g30145,g18386);
  OR2 OR2_1351(g24270,g23165,g18614);
  OR2 OR2_1352(g26911,g26612,g24230);
  OR4 OR4_48(I30741,g32085,g32030,g32224,g32013);
  OR2 OR2_1353(g30447,g29798,g21856);
  OR2 OR2_1354(g21894,g20112,g15107);
  OR2 OR2_1355(g34447,g34363,g18552);
  OR2 OR2_1356(g32995,g32330,g18375);
  OR2 OR2_1357(g24460,g10967,g22450);
  OR2 OR2_1358(g29904,g28312,g26146);
  OR2 OR2_1359(g13657,g7251,g10616);
  OR2 OR2_1360(g29252,g28712,g18486);
  OR2 OR2_1361(g28884,g27568,g16885);
  OR2 OR2_1362(g26785,g10776,g24468);
  OR2 OR2_1363(g24267,g23439,g18611);
  OR2 OR2_1364(g30451,g29877,g21860);
  OR2 OR2_1365(g30472,g30186,g21943);
  OR4 OR4_49(I30735,g32369,g32376,g32089,g32035);
  OR2 OR2_1366(g34629,g34495,g18654);
  OR4 OR4_50(g17569,g14416,g14394,g11995,I18492);
  OR2 OR2_1367(g34451,g34393,g18664);
  OR2 OR2_1368(g34628,g34493,g18653);
  OR2 OR2_1369(g34911,g34909,g18188);
  OR2 OR2_1370(g26950,g26357,g24288);
  OR2 OR2_1371(g22751,g19333,g15716);
  OR3 OR3_33(g27008,g26866,g21370,I25736);
  OR2 OR2_1372(g22639,g18950,g15612);
  OR2 OR2_1373(g27555,g26095,g24686);
  OR2 OR2_1374(g28580,g27328,g26275);
  OR2 OR2_1375(g29508,g28152,g27041);
  OR3 OR3_34(g8476,g1399,g1459,I12611);
  OR2 OR2_1376(g20160,g16163,g13415);
  OR2 OR2_1377(g30355,g30131,g18360);
  OR2 OR2_1378(g27570,g26126,g24722);
  OR2 OR2_1379(g31929,g31540,g22093);
  OR2 OR2_1380(g32989,g32241,g18326);
  OR2 OR2_1381(g30370,g30135,g18440);
  OR2 OR2_1382(g25629,g24962,g18258);
  OR2 OR2_1383(g27907,g17424,g26770);
  OR2 OR2_1384(g16959,g13542,g11142);
  OR2 OR2_1385(g31020,g29375,g28164);
  OR2 OR2_1386(g31928,g31517,g22092);
  OR2 OR2_1387(g14187,g8871,g11771);
  OR2 OR2_1388(g32988,g32232,g18325);
  OR2 OR2_1389(g28084,g27254,g18698);
  OR2 OR2_1390(g33020,g32160,g21734);
  OR2 OR2_1391(g33583,g33074,g18448);
  OR2 OR2_1392(g25628,g24600,g18249);
  OR2 OR2_1393(g25911,g22514,g24510);
  OR2 OR2_1394(g27239,g25881,g24465);
  OR2 OR2_1395(g19605,g15707,g13063);
  OR2 OR2_1396(g33046,g32308,g21912);
  OR2 OR2_1397(g32271,g31209,g29731);
  OR2 OR2_1398(g34172,g33795,g19914);
  OR4 OR4_51(g28179,g27494,g27474,g27445,g27421);
  OR2 OR2_1399(g27567,g26121,g24714);
  OR2 OR2_1400(g27238,g25879,g24464);
  OR4 OR4_52(g17510,g14393,g14362,g11972,I18449);
  OR2 OR2_1401(g30394,g29805,g21753);
  OR2 OR2_1402(g30367,g30133,g18418);
  OR2 OR2_1403(g24201,g22848,g18104);
  OR2 OR2_1404(g24277,g23188,g18647);
  OR2 OR2_1405(g25591,g24642,g21705);
  OR2 OR2_1406(g33282,g32143,g29577);
  OR4 OR4_53(g28186,g27209,g27185,g27161,g27146);
  OR2 OR2_1407(g28685,g27433,g16637);
  OR2 OR2_1408(g31302,g29590,g28302);
  OR2 OR2_1409(g28373,g27180,g15849);
  OR2 OR2_1410(g25754,g25179,g22101);
  OR2 OR2_1411(g30420,g29769,g21804);
  OR2 OR2_1412(g28417,g27219,g15881);
  OR2 OR2_1413(g24782,g23857,g23872);
  OR2 OR2_1414(g30446,g29788,g21855);
  OR2 OR2_1415(g34446,g34390,g18550);
  OR2 OR2_1416(g34318,g25850,g34063);
  OR2 OR2_1417(g28334,g27131,g15817);
  OR2 OR2_1418(g29756,g22717,g28223);
  OR2 OR2_1419(g24352,g22157,g18821);
  OR2 OR2_1420(g26902,g26378,g24219);
  OR2 OR2_1421(g26957,g26517,g24295);
  OR2 OR2_1422(g34025,g33927,g18672);
  OR2 OR2_1423(g31768,g30033,g30045);
  OR2 OR2_1424(g26377,g24700,g23007);
  OR2 OR2_1425(g30540,g30275,g22086);
  OR2 OR2_1426(g13295,g10625,g10655);
  OR2 OR2_1427(g15582,g8977,g12925);
  OR2 OR2_1428(g24266,g22329,g18561);
  OR2 OR2_1429(g32132,g31487,g31479);
  OR2 OR2_1430(g9535,g209,g538);
  OR2 OR2_1431(g31881,g31018,g21775);
  OR2 OR2_1432(g28216,g27036,g27043);
  OR2 OR2_1433(g24853,g21452,g24001);
  OR2 OR2_1434(g22684,g19206,g15703);
  OR2 OR2_1435(g32259,g31185,g29709);
  OR2 OR2_1436(g30377,g30124,g18472);
  OR2 OR2_1437(g32225,g30576,g29336);
  OR2 OR2_1438(g34957,g34948,g21662);
  OR2 OR2_1439(g34377,g26304,g34141);
  OR2 OR2_1440(g33027,g32314,g21796);
  OR3 OR3_35(I22912,g21555,g21364,g21357);
  OR2 OR2_1441(g31890,g31143,g21823);
  OR2 OR2_1442(g24401,g23811,g21298);
  OR2 OR2_1443(g30562,g30289,g22133);
  OR2 OR2_1444(g31249,g25971,g29523);
  OR2 OR2_1445(g19359,g17786,g14875);
  OR2 OR2_1446(g34645,g34556,g18786);
  OR2 OR2_1447(g19535,g15651,g13020);
  OR2 OR2_1448(g31248,g25970,g29522);
  OR2 OR2_1449(g28747,g27521,g13942);
  OR2 OR2_1450(g34290,g26848,g34219);
  OR2 OR2_1451(g33552,g33400,g18343);
  OR2 OR2_1452(g13289,g10619,g10624);
  OR2 OR2_1453(g33003,g32323,g18429);
  OR3 OR3_36(g33204,g32317,I30750,I30751);
  OR2 OR2_1454(g26895,g26783,g18148);
  OR2 OR2_1455(g31779,g30050,g28673);
  OR4 OR4_54(I31843,g33470,g33471,g33472,g33473);
  OR2 OR2_1456(g10800,g7517,g952);
  OR2 OR2_1457(g19344,g17771,g14832);
  OR2 OR2_1458(g27566,g26119,g24713);
  OR2 OR2_1459(g28814,g27545,g16841);
  OR2 OR2_1460(g30427,g29796,g21811);
  OR2 OR2_1461(g20276,g16243,g13566);
  OR2 OR2_1462(g29583,g28182,g27099);
  OR2 OR2_1463(g32375,g29896,g31324);
  OR2 OR2_1464(g14936,g10776,g8703);
  OR2 OR2_1465(g30366,g30122,g18417);
  OR4 OR4_55(I30054,g29385,g31376,g30735,g30825);
  OR2 OR2_1466(g24276,g23083,g18646);
  OR2 OR2_1467(g28751,g27526,g16766);
  OR2 OR2_1468(g28772,g27534,g16802);
  OR2 OR2_1469(g34366,g26257,g34133);
  OR4 OR4_56(I31869,g33519,g33520,g33521,g33522);
  OR2 OR2_1470(g34632,g34565,g15119);
  OR2 OR2_1471(g25739,g25149,g22054);
  OR2 OR2_1472(g24254,g23265,g18306);
  OR4 OR4_57(I31868,g33515,g33516,g33517,g33518);
  OR2 OR2_1473(g28230,g27669,g14261);
  OR2 OR2_1474(g33945,g32430,g33455);
  OR2 OR2_1475(g25738,g25059,g22053);
  OR2 OR2_1476(g25645,g24679,g21738);
  OR2 OR2_1477(g30547,g30194,g22118);
  OR2 OR2_1478(g30403,g29750,g21762);
  OR2 OR2_1479(g33999,g33893,g18436);
  OR2 OR2_1480(g33380,g32234,g29926);
  OR2 OR2_1481(g25699,g25125,g21918);
  OR2 OR2_1482(g34403,g34180,g25085);
  OR2 OR2_1483(g29282,g28617,g18745);
  OR2 OR2_1484(g28416,g27218,g15880);
  OR2 OR2_1485(g16261,g7898,g13469);
  OR2 OR2_1486(g32994,g32290,g18367);
  OR2 OR2_1487(g33998,g33878,g18428);
  OR2 OR2_1488(g29302,g28601,g18798);
  OR2 OR2_1489(g25698,g25104,g21917);
  OR2 OR2_1490(g29105,g27645,g17134);
  OR2 OR2_1491(g30481,g30221,g21977);
  OR2 OR2_1492(g7932,g4072,g4153);
  OR2 OR2_1493(g26956,g26487,g24294);
  OR2 OR2_1494(g30551,g30235,g22122);
  OR4 OR4_58(I30734,g31790,g32191,g32086,g32095);
  OR2 OR2_1495(g26889,g26689,g24195);
  OR2 OR2_1496(g31932,g31792,g22107);
  OR2 OR2_1497(g26888,g26671,g24194);
  OR3 OR3_37(g23721,g21401,g21385,I22852);
  OR2 OR2_1498(g25632,g24558,g18277);
  OR2 OR2_1499(g28578,g27327,g26273);
  OR2 OR2_1500(g30127,g28494,g16805);
  OR2 OR2_1501(g29768,g22760,g28229);
  OR2 OR2_1502(g34127,g33657,g32438);
  OR2 OR2_1503(g31897,g31237,g24322);
  OR2 OR2_1504(g30490,g30167,g21986);
  OR2 OR2_1505(g33961,g33789,g21712);
  OR2 OR2_1506(g25661,g24754,g21786);
  OR2 OR2_1507(g27484,g25988,g24628);
  OR2 OR2_1508(g30376,g30112,g18471);
  OR2 OR2_1509(g30385,g30172,g18518);
  OR2 OR2_1510(g26931,g26778,g18547);
  OR2 OR2_1511(g30103,g28477,g16731);
  OR2 OR2_1512(g34376,g26301,g34140);
  OR2 OR2_1513(g34297,g26858,g34228);
  OR2 OR2_1514(g34103,g33701,g33707);
  OR2 OR2_1515(g33026,g32307,g21795);
  OR2 OR2_1516(g30354,g30064,g18359);
  OR2 OR2_1517(g22516,g21559,g12817);
  OR2 OR2_1518(g34980,g34969,g18587);
  OR3 OR3_38(g33212,g32328,I30755,I30756);
  OR2 OR2_1519(g25715,g25071,g21966);
  OR2 OR2_1520(g8679,g222,g199);
  OR2 OR2_1521(g34095,g33681,g33687);
  OR2 OR2_1522(g30824,g13833,g29789);
  OR2 OR2_1523(g28720,g27486,g16704);
  OR2 OR2_1524(g28041,g24145,g26878);
  OR2 OR2_1525(g17264,g7118,g14309);
  OR2 OR2_1526(g28430,g27229,g15914);
  OR2 OR2_1527(g32125,g30918,g29376);
  OR2 OR2_1528(g28746,g27520,g16762);
  OR2 OR2_1529(g32977,g32169,g21710);
  OR2 OR2_1530(g19604,g15704,g13059);
  OR4 OR4_59(I30469,g31672,g31710,g31021,g30937);
  OR2 OR2_1531(g29249,g28658,g18438);
  OR2 OR2_1532(g26089,g24501,g22534);
  OR2 OR2_1533(g24907,g21558,g24015);
  OR4 OR4_60(I30468,g29385,g31376,g30735,g30825);
  OR2 OR2_1534(g29482,g28524,g27588);
  OR2 OR2_1535(g34931,g2984,g34912);
  OR2 OR2_1536(g29248,g28677,g18434);
  OR3 OR3_39(g33149,g32204,I30717,I30718);
  OR2 OR2_1537(g30426,g29785,g21810);
  OR2 OR2_1538(g32353,g29853,g31283);
  OR2 OR2_1539(g33387,g32263,g29954);
  OR2 OR2_1540(g24239,g22752,g18250);
  OR2 OR2_1541(g9055,g2606,g2625);
  OR2 OR2_1542(g28684,g27432,g16636);
  OR2 OR2_1543(g32144,g30927,g30930);
  OR2 OR2_1544(g33620,g33360,g18774);
  OR2 OR2_1545(g34190,g33802,g33810);
  OR2 OR2_1546(g24238,g23254,g18248);
  OR2 OR2_1547(g30520,g30272,g22041);
  OR2 OR2_1548(g28517,g27280,g26154);
  OR2 OR2_1549(g30546,g30277,g22117);
  OR2 OR2_1550(g33971,g33890,g18330);
  OR2 OR2_1551(g29786,g22843,g28240);
  OR2 OR2_1552(g25671,g24637,g21828);
  OR2 OR2_1553(g34024,g33807,g24331);
  OR2 OR2_1554(g13938,g11213,g11191);
  OR2 OR2_1555(g24518,g22517,g7601);
  OR2 OR2_1556(g22530,g16751,g20171);
  OR2 OR2_1557(g28362,g27154,g15840);
  OR2 OR2_1558(g30497,g30242,g21993);
  OR2 OR2_1559(g24935,g22937,g19749);
  OR4 OR4_61(I12903,g4222,g4219,g4216,g4213);
  OR2 OR2_1560(g29233,g28171,g18234);
  OR2 OR2_1561(g26969,g26313,g24329);
  OR3 OR3_40(I18421,g14447,g14417,g14395);
  OR2 OR2_1562(g32289,g24796,g31230);
  OR2 OR2_1563(g22641,g18974,g15631);
  OR2 OR2_1564(g34625,g34532,g18610);
  OR2 OR2_1565(g26968,g26307,g24321);
  OR4 OR4_62(g17464,g14334,g14313,g11935,I18385);
  OR2 OR2_1566(g31896,g31242,g24305);
  OR2 OR2_1567(g34250,g34111,g21713);
  OR2 OR2_1568(g32288,g31226,g31229);
  OR2 OR2_1569(g28727,g27500,g16729);
  OR2 OR2_1570(g16258,g13247,g10856);
  OR2 OR2_1571(g33011,g32338,g18481);
  OR2 OR2_1572(g30339,g29629,g18244);
  OR2 OR2_1573(g24215,g23484,g18196);
  OR2 OR2_1574(g24577,g2856,g22531);
  OR2 OR2_1575(g30338,g29613,g18240);
  OR2 OR2_1576(g34644,g34555,g18769);
  OR2 OR2_1577(g33582,g33351,g18444);
  OR2 OR2_1578(g19534,g15650,g13019);
  OR2 OR2_1579(g27241,g24584,g25984);
  OR2 OR2_1580(g28347,g27138,g15822);
  OR2 OR2_1581(g29717,g28200,g10883);
  OR2 OR2_1582(g33310,g29631,g32165);
  OR2 OR2_1583(g26894,g25979,g18129);
  OR2 OR2_1584(g33627,g33376,g18826);
  OR2 OR2_1585(g31925,g31789,g22061);
  OR2 OR2_1586(g32976,g32207,g21704);
  OR2 OR2_1587(g32985,g31963,g18266);
  OR2 OR2_1588(g24349,g23646,g18805);
  OR2 OR2_1589(g16810,g13461,g11032);
  OR2 OR2_1590(g25700,g25040,g21919);
  OR2 OR2_1591(g28600,g27339,g16427);
  OR2 OR2_1592(g25659,g24707,g21784);
  OR2 OR2_1593(g25625,g24553,g18226);
  OR2 OR2_1594(g20083,g2902,g17058);
  OR2 OR2_1595(g30527,g30192,g22073);
  OR2 OR2_1596(g30411,g29872,g21770);
  OR2 OR2_1597(g33050,g31974,g21930);
  OR2 OR2_1598(g32374,g29895,g31323);
  OR3 OR3_41(g33958,g33532,I31873,I31874);
  OR2 OR2_1599(g24348,g22149,g18804);
  OR2 OR2_1600(g34411,g34186,g25142);
  OR2 OR2_1601(g16970,g13567,g11163);
  OR2 OR2_1602(g25658,g24635,g21783);
  OR2 OR2_1603(g28372,g27178,g15848);
  OR2 OR2_1604(g23217,g19588,g16023);
  OR2 OR2_1605(g33386,g32258,g29951);
  OR2 OR2_1606(g26910,g26571,g24228);
  OR2 OR2_1607(g33603,g33372,g18515);
  OR2 OR2_1608(g25943,g24423,g22299);
  OR4 OR4_63(I30740,g31776,g32188,g32083,g32087);
  OR2 OR2_1609(g13623,g482,g12527);
  OR2 OR2_1610(g25644,g24622,g21737);
  OR2 OR2_1611(g30503,g30243,g22024);
  OR2 OR2_1612(g28063,g27541,g21773);
  OR2 OR2_1613(g34894,g34862,g21678);
  OR2 OR2_1614(g29148,g27651,g26606);
  OR2 OR2_1615(g32392,g31513,g30000);
  OR2 OR2_1616(g27515,g26051,g13431);
  OR2 OR2_1617(g30450,g29861,g21859);
  OR2 OR2_1618(g24653,g2848,g22585);
  OR2 OR2_1619(g34450,g34281,g18663);
  OR2 OR2_1620(g13155,g11496,g11546);
  OR2 OR2_1621(g31793,g28031,g30317);
  OR2 OR2_1622(g34819,g34741,g34684);
  OR2 OR2_1623(g34257,g34226,g18674);
  OR2 OR2_1624(g28209,g27223,g27141);
  OR2 OR2_1625(g30496,g30231,g21992);
  OR2 OR2_1626(g8956,g1913,g1932);
  OR2 OR2_1627(g34979,g34875,g34968);
  OR2 OR2_1628(g34055,g33909,g33910);
  OR2 OR2_1629(g33549,g33328,g18337);
  OR2 OR2_1630(g28208,g27025,g27028);
  OR2 OR2_1631(g26877,g21658,g25577);
  OR2 OR2_1632(g34978,g34874,g34967);
  OR2 OR2_1633(g33548,g33327,g18336);
  OR2 OR2_1634(g27584,g26165,g24758);
  OR2 OR2_1635(g25867,g25449,g23884);
  OR2 OR2_1636(g25894,g24817,g23229);
  OR2 OR2_1637(g30384,g30101,g18517);
  OR2 OR2_1638(g31317,g29611,g29626);
  OR2 OR2_1639(g33317,g29688,g32179);
  OR2 OR2_1640(g29229,g28532,g18191);
  OR2 OR2_1641(g25714,g25056,g21965);
  OR2 OR2_1642(g28614,g27351,g26311);
  OR2 OR2_1643(g25707,g25041,g18749);
  OR2 OR2_1644(g25819,g25323,g23836);
  OR2 OR2_1645(g28607,g27342,g26303);
  OR2 OR2_1646(g29228,g28426,g18173);
  OR2 OR2_1647(g25910,g25565,g22142);
  OR2 OR2_1648(g28320,g27116,g15808);
  OR2 OR2_1649(g31002,g29362,g28154);
  OR2 OR2_1650(g28073,g27097,g21875);
  OR2 OR2_1651(g33002,g32304,g18419);
  OR2 OR2_1652(g33057,g31968,g22019);
  OR2 OR2_1653(g34801,g34756,g18588);
  OR2 OR2_1654(g34735,g34709,g15116);
  OR2 OR2_1655(g32124,g24488,g30920);
  OR2 OR2_1656(g29716,g28199,g15856);
  OR2 OR2_1657(g24200,g22831,g18103);
  OR2 OR2_1658(g31245,g25964,g29516);
  OR2 OR2_1659(g34019,g33889,g18506);
  OR2 OR2_1660(g26917,g26122,g18233);
  OR2 OR2_1661(g15792,g12920,g10501);
  OR3 OR3_42(g26866,g20204,g20242,g24363);
  OR2 OR2_1662(g28565,g27315,g26253);
  OR2 OR2_1663(g33626,g33374,g18825);
  OR2 OR2_1664(g33323,g31936,g32442);
  OR2 OR2_1665(g34695,g34523,g34322);
  OR2 OR2_1666(g25590,g21694,g24160);
  OR2 OR2_1667(g34018,g33887,g18505);
  OR2 OR2_1668(g30526,g30181,g22072);
  OR2 OR2_1669(g32267,g31208,g31218);
  OR2 OR2_1670(g32294,g31231,g31232);
  OR2 OR2_1671(g33298,g32158,g29622);
  OR2 OR2_1672(g25741,g25178,g22056);
  OR2 OR2_1673(g28641,g27385,g16591);
  OR2 OR2_1674(g31775,g30048,g30059);
  OR4 OR4_64(I30123,g29385,g31376,g30735,g30825);
  OR2 OR2_1675(g8957,g2338,g2357);
  OR2 OR2_1676(g24799,g23901,g23921);
  OR2 OR2_1677(g30402,g29871,g21761);
  OR2 OR2_1678(g24813,g22685,g19594);
  OR4 OR4_65(I30751,g32042,g32161,g31943,g31959);
  OR2 OR2_1679(g30457,g29369,g21885);
  OR2 OR2_1680(g34402,g34179,g25084);
  OR2 OR2_1681(g34457,g34394,g18670);
  OR2 OR2_1682(g26923,g25923,g18290);
  OR2 OR2_1683(g32219,g31131,g29620);
  OR2 OR2_1684(g33232,g32034,g30936);
  OR2 OR2_1685(g25735,g25077,g18783);
  OR2 OR2_1686(g25877,g25502,g23919);
  OR2 OR2_1687(g28635,g27375,g16537);
  OR2 OR2_1688(g32218,g31130,g29619);
  OR2 OR2_1689(g27135,g24387,g25803);
  OR2 OR2_1690(g33995,g33848,g18425);
  OR2 OR2_1691(g34001,g33844,g18450);
  OR2 OR2_1692(g33261,g32111,g29525);
  OR2 OR2_1693(g25695,g24998,g21914);
  OR2 OR2_1694(g31880,g31280,g21774);
  OR2 OR2_1695(g30597,g13564,g29693);
  OR2 OR2_1696(g34256,g34173,g24303);
  OR2 OR2_1697(g29802,g28243,g22871);
  OR2 OR2_1698(g34280,g26833,g34213);
  OR2 OR2_1699(g29730,g28150,g28141);
  OR2 OR2_1700(g30300,g28246,g27252);
  OR2 OR2_1701(g29793,g28237,g27247);
  OR2 OR2_1702(g34624,g34509,g18592);
  OR2 OR2_1703(g34300,g26864,g34230);
  OR2 OR2_1704(g15125,g10363,g13605);
  OR2 OR2_1705(g26876,g21655,g25576);
  OR2 OR2_1706(g26885,g26541,g24191);
  OR3 OR3_43(g23751,g21415,g21402,I22880);
  OR2 OR2_1707(g25917,g22524,g24518);
  OR2 OR2_1708(g32277,g31211,g29733);
  OR2 OR2_1709(g24214,g23471,g18195);
  OR2 OR2_1710(g31316,g29609,g29624);
  OR2 OR2_1711(g33316,g29685,g32178);
  OR2 OR2_1712(g22634,g18934,g15590);
  OR2 OR2_1713(g24207,g23396,g18119);
  OR2 OR2_1714(g22872,g19372,g19383);
  OR4 OR4_66(I29985,g29385,g31376,g30735,g30825);
  OR3 OR3_44(I22958,g21603,g21386,g21365);
  OR2 OR2_1715(g34231,g33898,g33902);
  OR2 OR2_1716(g29504,g28143,g25875);
  OR2 OR2_1717(g25706,g25030,g18748);
  OR2 OR2_1718(g25597,g24892,g21719);
  OR2 OR2_1719(g32037,g30566,g29329);
  OR2 OR2_1720(g33989,g33870,g18398);
  OR2 OR2_1721(g33056,g32327,g22004);
  OR2 OR2_1722(g13570,g9223,g11130);
  OR2 OR2_1723(g25689,g24849,g21888);
  OR2 OR2_1724(g13914,g8643,g11380);
  OR2 OR2_1725(g33611,g33243,g18632);
  OR2 OR2_1726(g31924,g31486,g22049);
  OR2 OR2_1727(g32984,g31934,g18264);
  OR2 OR2_1728(g33988,g33861,g18397);
  OR2 OR2_1729(g25688,g24812,g21887);
  OR2 OR2_1730(g28750,g27525,g16765);
  OR2 OR2_1731(g25624,g24408,g18224);
  OR2 OR2_1732(g26916,g25916,g18232);
  OR2 OR2_1733(g30511,g30180,g22032);
  OR2 OR2_1734(g20241,g16233,g13541);
  OR2 OR2_1735(g32352,g29852,g31282);
  OR4 OR4_67(I30746,g32047,g31985,g31991,g32309);
  OR2 OR2_1736(g24241,g22920,g18252);
  OR2 OR2_1737(g33271,g32120,g29549);
  OR2 OR2_1738(g27972,g26131,g26105);
  OR2 OR2_1739(g32155,g30935,g29475);
  OR2 OR2_1740(g15017,g10776,g8703);
  OR2 OR2_1741(g28091,g27665,g21913);
  OR2 OR2_1742(g32266,g30604,g29354);
  OR2 OR2_1743(g29245,g28676,g18384);
  OR2 OR2_1744(g26721,g10776,g24444);
  OR2 OR2_1745(g29299,g28587,g18794);
  OR2 OR2_1746(g33031,g32315,g21841);
  OR2 OR2_1747(g30456,g29378,g21869);
  OR2 OR2_1748(g34456,g34395,g18669);
  OR2 OR2_1749(g29298,g28571,g18793);
  OR2 OR2_1750(g24235,g22632,g18238);
  OR2 OR2_1751(g13941,g11019,g11023);
  OR2 OR2_1752(g31887,g31292,g21820);
  OR2 OR2_1753(g28390,g27207,g15861);
  OR2 OR2_1754(g30480,g29321,g21972);
  OR2 OR2_1755(g30916,g13853,g29799);
  OR2 OR2_1756(g29775,g25966,g28232);
  OR4 OR4_68(I26523,g20720,g20857,g20998,g21143);
  OR2 OR2_1757(g25885,g25522,g23957);
  OR2 OR2_1758(g30550,g30226,g22121);
  OR2 OR2_1759(g30314,g28268,g27266);
  OR2 OR2_1760(g23615,g20109,g20131);
  OR2 OR2_1761(g30287,g28653,g27677);
  OR2 OR2_1762(g34314,g25831,g34061);
  OR2 OR2_1763(g30307,g28256,g27260);
  OR2 OR2_1764(g33393,g32286,g29984);
  OR2 OR2_1765(g23720,g20165,g16801);
  OR4 OR4_69(I12902,g4235,g4232,g4229,g4226);
  OR2 OR2_1766(g25763,g25113,g18817);
  OR2 OR2_1767(g29232,g28183,g18231);
  OR2 OR2_1768(g31764,g30015,g30032);
  OR2 OR2_1769(g23275,g19680,g16160);
  OR2 OR2_1770(g34721,g34696,g18135);
  OR2 OR2_1771(g31869,g30592,g18221);
  OR4 OR4_70(I30193,g31070,g30614,g30673,g31528);
  OR2 OR2_1772(g30431,g29875,g21815);
  OR2 OR2_1773(g33960,g33759,g21701);
  OR2 OR2_1774(g25660,g24726,g21785);
  OR2 OR2_1775(g29261,g28247,g18605);
  OR2 OR2_1776(g31868,g30600,g18204);
  OR2 OR2_1777(g26335,g1526,g24609);
  OR2 OR2_1778(g19572,g17133,g14193);
  OR2 OR2_1779(g22152,g21188,g17469);
  OR2 OR2_1780(g26930,g26799,g18544);
  OR2 OR2_1781(g34269,g34083,g18732);
  OR2 OR2_1782(g30341,g29380,g18246);
  OR2 OR2_1783(g26694,g24444,g10704);
  OR2 OR2_1784(g26965,g26336,g24317);
  OR2 OR2_1785(g33709,g32414,g33441);
  OR2 OR2_1786(g34268,g34082,g18730);
  OR2 OR2_1787(g31259,g25992,g29554);
  OR2 OR2_1788(g32285,g31222,g29740);
  OR2 OR2_1789(g33259,g32109,g29521);
  OR2 OR2_1790(g28536,g27293,g26205);
  OR4 OR4_71(I30727,g31759,g32196,g31933,g31941);
  OR2 OR2_1791(g31258,g25991,g29550);
  OR2 OR2_1792(g24206,g23386,g18110);
  OR2 OR2_1793(g13728,g6804,g12527);
  OR2 OR2_1794(g28702,g27457,g16670);
  OR2 OR2_1795(g30734,g13808,g29774);
  OR3 OR3_45(I22298,g20371,g20161,g20151);
  OR2 OR2_1796(g30335,g29746,g18174);
  OR2 OR2_1797(g34734,g34681,g18652);
  OR2 OR2_1798(g25721,g25057,g18766);
  OR2 OR2_1799(g28621,g27359,g16518);
  OR2 OR2_1800(g25596,g24865,g21718);
  OR4 OR4_72(I31853,g33488,g33489,g33490,g33491);
  OR2 OR2_1801(g33043,g32195,g24325);
  OR2 OR2_1802(g31244,g25963,g29515);
  OR2 OR2_1803(g20082,g16026,g13321);
  OR2 OR2_1804(g28564,g27314,g26252);
  OR2 OR2_1805(g23193,g19556,g15937);
  OR4 OR4_73(I23756,g23457,g23480,g23494,g23511);
  OR2 OR2_1806(g26278,g24545,g24549);
  OR2 OR2_1807(g33069,g32009,g22113);
  OR2 OR2_1808(g33602,g33425,g18511);
  OR2 OR2_1809(g25942,g24422,g22298);
  OR2 OR2_1810(g31774,g30046,g30057);
  OR2 OR2_1811(g7834,g2886,g2946);
  OR2 OR2_1812(g30487,g30187,g21983);
  OR2 OR2_1813(g31375,g29628,g28339);
  OR2 OR2_1814(g33068,g31994,g22112);
  OR3 OR3_46(g33955,g33505,I31858,I31859);
  OR2 OR2_1815(g24345,g23606,g18788);
  OR2 OR2_1816(g25655,g24645,g18607);
  OR2 OR2_1817(g31879,g31475,g21745);
  OR2 OR2_1818(g30502,g30232,g22023);
  OR2 OR2_1819(g28062,g27288,g21746);
  OR2 OR2_1820(g30557,g30247,g22128);
  OR2 OR2_1821(g33970,g33868,g18322);
  OR2 OR2_1822(g34619,g34528,g18581);
  OR3 OR3_47(I22880,g21509,g21356,g21351);
  OR2 OR2_1823(g25670,g24967,g18626);
  OR2 OR2_1824(g29271,g28333,g18637);
  OR2 OR2_1825(g31878,g31015,g21733);
  OR4 OR4_74(I31864,g33510,g33511,g33512,g33513);
  OR2 OR2_1826(g30443,g29808,g21852);
  OR2 OR2_1827(g34618,g34527,g18580);
  OR2 OR2_1828(g24398,g23801,g21296);
  OR2 OR2_1829(g30279,g28637,g27668);
  OR2 OR2_1830(g34443,g34385,g18545);
  OR2 OR2_1831(g25734,g25058,g18782);
  OR2 OR2_1832(g28634,g27374,g16536);
  OR2 OR2_1833(g28851,g27558,g16870);
  OR2 OR2_1834(g31886,g31481,g21791);
  OR2 OR2_1835(g29753,g28213,g22720);
  OR4 OR4_75(g25839,g25507,g25485,g25459,g25420);
  OR2 OR2_1836(g34278,g26829,g34212);
  OR2 OR2_1837(g30469,g30153,g21940);
  OR2 OR2_1838(g33967,g33842,g18319);
  OR2 OR2_1839(g33994,g33841,g18424);
  OR2 OR2_1840(g27506,g26021,g24639);
  OR2 OR2_1841(g30286,g28191,g28186);
  OR2 OR2_1842(g25694,g24638,g18738);
  OR2 OR2_1843(g25667,g24682,g18619);
  OR2 OR2_1844(g24263,g23497,g18529);
  OR2 OR2_1845(g34286,g26842,g34216);
  OR2 OR2_1846(g30468,g30238,g21939);
  OR2 OR2_1847(g34468,g34342,g18718);
  OR2 OR2_1848(g34039,g33743,g18736);
  OR2 OR2_1849(g34306,g25782,g34054);
  OR4 OR4_76(g29529,g28303,g28293,g28283,g28267);
  OR2 OR2_1850(g22640,g18951,g15613);
  OR2 OR2_1851(g34038,g33731,g18735);
  OR2 OR2_1852(g31919,g31758,g22044);
  OR2 OR2_1853(g32454,g30322,g31795);
  OR2 OR2_1854(g25619,g24961,g18193);
  OR2 OR2_1855(g15124,g13605,g4581);
  OR2 OR2_1856(g26884,g26511,g24190);
  OR2 OR2_1857(g28574,g27324,g26270);
  OR2 OR2_1858(g31918,g31786,g22015);
  OR2 OR2_1859(g28047,g27676,g18160);
  OR2 OR2_1860(g33010,g32301,g18473);
  OR2 OR2_1861(g34601,g34488,g18211);
  OR2 OR2_1862(g29764,g28219,g28226);
  OR2 OR2_1863(g25618,g25491,g18192);
  OR2 OR2_1864(g34975,g34871,g34964);
  OR2 OR2_1865(g24500,g24011,g21605);
  OR2 OR2_1866(g33545,g33399,g18324);
  OR2 OR2_1867(g9013,g2472,g2491);
  OR2 OR2_1868(g26363,g2965,g24965);
  OR2 OR2_1869(g33599,g33087,g18500);
  OR2 OR2_1870(g32239,g30595,g29350);
  OR2 OR2_1871(g28051,g27699,g18166);
  OR2 OR2_1872(g27240,g25883,g24467);
  OR2 OR2_1873(g28072,g27086,g21874);
  OR2 OR2_1874(g33598,g33364,g18496);
  OR2 OR2_1875(g32238,g30594,g29349);
  OR4 OR4_77(I29352,g29322,g29315,g30315,g30308);
  OR2 OR2_1876(g28592,g27333,g26288);
  OR4 OR4_78(I31874,g33528,g33529,g33530,g33531);
  OR2 OR2_1877(g34791,g34771,g18184);
  OR2 OR2_1878(g22662,g19069,g15679);
  OR2 OR2_1879(g34884,g34858,g21666);
  OR2 OR2_1880(g29259,g28304,g18603);
  OR2 OR2_1881(g29225,g28451,g18158);
  OR2 OR2_1882(g30410,g29857,g21769);
  OR2 OR2_1883(g31322,g26128,g29635);
  OR2 OR2_1884(g14062,g11047,g11116);
  OR2 OR2_1885(g34168,g33787,g19784);
  OR2 OR2_1886(g27563,g26104,g24704);
  OR2 OR2_1887(g29258,g28238,g18601);
  OR2 OR2_1888(g31901,g31516,g21909);
  OR2 OR2_1889(g33159,g32016,g30730);
  OR2 OR2_1890(g30479,g29320,g21950);
  OR2 OR2_1891(g33977,g33876,g18348);
  OR2 OR2_1892(g30363,g30121,g18407);
  OR2 OR2_1893(g25601,g24660,g18112);
  OR2 OR2_1894(g12981,g12219,g9967);
  OR2 OR2_1895(g24273,g23166,g18630);
  OR2 OR2_1896(g25677,g24684,g21834);
  OR2 OR2_1897(g31783,I29351,I29352);
  OR2 OR2_1898(g23209,g19585,g19601);
  OR2 OR2_1899(g30478,g30248,g21949);
  OR2 OR2_1900(g34015,g33858,g18502);
  OR2 OR2_1901(g29244,g28692,g18380);
  OR2 OR2_1902(g33561,g33408,g18376);
  OR2 OR2_1903(g30486,g30177,g21982);
  OR2 OR2_1904(g31295,g26090,g29598);
  OR2 OR2_1905(g26922,g25902,g18288);
  OR2 OR2_1906(g28731,g27504,g16733);
  OR2 OR2_1907(g33295,g32153,g29605);
  OR2 OR2_1908(g31144,g29477,g28193);
  OR2 OR2_1909(g25937,g24406,g22216);
  OR2 OR2_1910(g30556,g30236,g22127);
  OR2 OR2_1911(g24234,g22622,g18237);
  OR2 OR2_1912(g13973,g11024,g11028);
  OR2 OR2_1913(g29068,g27628,g17119);
  OR4 OR4_79(g25791,g25411,g25371,g25328,g25290);
  OR2 OR2_1914(g28691,g27437,g16642);
  OR2 OR2_1915(g29879,g28289,g26096);
  OR2 OR2_1916(g26953,g26486,g24291);
  OR2 OR2_1917(g28405,g27216,g15875);
  OR2 OR2_1918(g33966,g33837,g18318);
  OR2 OR2_1919(g25666,g24788,g21793);
  OR2 OR2_1920(g33017,g32292,g18510);
  OR2 OR2_1921(g26800,g24922,g24929);
  OR2 OR2_1922(g34321,g25866,g34065);
  OR2 OR2_1923(g30531,g30274,g22077);
  OR2 OR2_1924(g23346,g19736,g16204);
  OR2 OR2_1925(g29792,g28235,g28244);
  OR2 OR2_1926(g12832,g10347,g10348);
  OR2 OR2_1927(g13761,g490,g12527);
  OR2 OR2_1928(g16022,g13048,g10707);
  OR2 OR2_1929(g26334,g1171,g24591);
  OR2 OR2_1930(g28046,g27667,g18157);
  OR2 OR2_1931(g32349,g29840,g31275);
  OR2 OR2_1932(g31289,g29580,g29591);
  OR2 OR2_1933(g30373,g30111,g18461);
  OR2 OR2_1934(g33289,g32148,g29588);
  OR2 OR2_1935(g22331,g21405,g17809);
  OR2 OR2_1936(g26964,g26259,g24316);
  OR2 OR2_1937(g34373,g26292,g34138);
  OR2 OR2_1938(g33023,g32313,g21751);
  OR2 OR2_1939(g31288,g2955,g29914);
  OR2 OR2_1940(g23153,g19521,g15876);
  OR2 OR2_1941(g33288,g32147,g29587);
  OR2 OR2_1942(g31308,g26101,g29614);
  OR2 OR2_1943(g33571,g33367,g18409);
  OR2 OR2_1944(g30417,g29874,g21801);
  OR2 OR2_1945(g34800,g34752,g18586);
  OR2 OR2_1946(g34417,g27678,g34196);
  OR2 OR2_1947(g28357,g27148,g15836);
  OR2 OR2_1948(g30334,g29837,g18143);
  OR2 OR2_1949(g28105,g27997,g22135);
  OR2 OR2_1950(g28743,g27517,g16758);
  OR2 OR2_1951(g29078,g27633,g26572);
  OR2 OR2_1952(g26909,g26543,g24227);
  OR3 OR3_48(I18385,g14413,g14391,g14360);
  OR2 OR2_1953(g34762,g34687,g34524);
  OR2 OR2_1954(g25740,g25164,g22055);
  OR2 OR2_1955(g26908,g26358,g24225);
  OR2 OR2_1956(g28640,g27384,g16590);
  OR2 OR2_1957(g30423,g29887,g21807);
  OR2 OR2_1958(g33976,g33869,g18347);
  OR2 OR2_1959(g33985,g33896,g18382);
  OR3 OR3_49(g24946,g22360,g22409,g8130);
  OR2 OR2_1960(g25676,g24668,g21833);
  OR2 OR2_1961(g25685,g24476,g21866);
  OR4 OR4_80(I30750,g31788,g32310,g32054,g32070);
  OR3 OR3_50(g33954,g33496,I31853,I31854);
  OR2 OR2_1962(g21891,g19948,g15103);
  OR2 OR2_1963(g24344,g22145,g18787);
  OR2 OR2_1964(g25654,g24634,g18606);
  OR2 OR2_1965(g25936,g24403,g22209);
  OR2 OR2_1966(g30543,g29338,g22110);
  OR4 OR4_81(I26522,g19890,g19935,g19984,g26365);
  OR2 OR2_1967(g31260,g25993,g29555);
  OR2 OR2_1968(g34000,g33943,g18441);
  OR2 OR2_1969(g26751,g24903,g24912);
  OR2 OR2_1970(g33260,g32110,g29524);
  OR2 OR2_1971(g29295,g28663,g18780);
  OR2 OR2_1972(g31668,g29924,g28558);
  OR2 OR2_1973(g14583,g10685,g542);
  OR2 OR2_1974(g25762,g25095,g18816);
  OR2 OR2_1975(g28662,g27407,g16612);
  OR2 OR2_1976(g26293,g24550,g24555);
  OR2 OR2_1977(g33559,g33073,g18368);
  OR4 OR4_82(I30192,g29385,g31376,g30735,g30825);
  OR2 OR2_1978(g33016,g32284,g18509);
  OR2 OR2_1979(g25587,g21682,g24157);
  OR2 OR2_1980(g33558,g33350,g18364);
  OR2 OR2_1981(g23750,g20174,g16840);
  OR2 OR2_1982(g31893,g31490,g21837);
  OR2 OR2_1983(g34807,g34764,g18596);
  OR2 OR2_1984(g34974,g34870,g34963);
  OR2 OR2_1985(g31865,g31149,g21709);
  OR2 OR2_1986(g33544,g33392,g18317);
  OR2 OR2_1987(g34639,g34486,g18722);
  OR2 OR2_1988(g12911,g10278,g12768);
  OR2 OR2_1989(g30293,g28236,g27246);
  OR3 OR3_51(g23796,g21462,g21433,I22958);
  OR2 OR2_1990(g28778,g27540,g16808);
  OR2 OR2_1991(g16239,g7892,g13432);
  OR2 OR2_1992(g34293,g26854,g34224);
  OR2 OR2_1993(g34638,g34484,g18721);
  OR2 OR2_1994(g34265,g34117,g18711);
  OR2 OR2_1995(g30416,g29858,g21800);
  OR2 OR2_1996(g27591,g26181,g24765);
  OR2 OR2_1997(g34416,g34191,g25159);
  OR2 OR2_1998(g29289,g28642,g18763);
  OR2 OR2_1999(g25747,g25130,g18795);
  OR2 OR2_2000(g28647,g27389,g16596);
  OR2 OR2_2001(g33610,g33242,g18616);
  OR2 OR2_2002(g29309,g28722,g18818);
  OR2 OR2_2003(g30391,g30080,g18557);
  OR2 OR2_2004(g33042,g32193,g24324);
  OR2 OR2_2005(g27147,g25802,g24399);
  OR2 OR2_2006(g31255,g25982,g29536);
  OR2 OR2_2007(g29288,g28630,g18762);
  OR2 OR2_2008(g33255,g32106,g29514);
  OR2 OR2_2009(g29224,g28919,g18156);
  OR2 OR2_2010(g30510,g30263,g22031);
  OR2 OR2_2011(g29308,g28612,g18815);
  OR2 OR2_2012(g24240,g22861,g18251);
  OR2 OR2_2013(g33270,g32119,g29547);
  OR2 OR2_2014(g28090,g27275,g18733);
  OR2 OR2_2015(g30579,g30173,g14571);
  OR2 OR2_2016(g27858,g17405,g26737);
  OR2 OR2_2017(g25751,g25061,g22098);
  OR2 OR2_2018(g28651,g27392,g16599);
  OR2 OR2_2019(g29495,g28563,g27614);
  OR2 OR2_2020(g33383,g32244,g29940);
  OR2 OR2_2021(g25639,g25122,g18530);
  OR2 OR2_2022(g34014,g33647,g18493);
  OR2 OR2_2023(g33030,g32166,g21826);
  OR2 OR2_2024(g31267,g29548,g28263);
  OR2 OR2_2025(g25638,g24977,g18316);
  OR2 OR2_2026(g34007,g33640,g18467);
  OR2 OR2_2027(g16883,g13509,g11115);
  OR2 OR2_2028(g33267,g32115,g29535);
  OR2 OR2_2029(g33294,g32152,g29604);
  OR2 OR2_2030(g27394,g25957,g24573);
  OR2 OR2_2031(g28331,g27129,g15814);
  OR2 OR2_2032(g30442,g29797,g21851);
  OR2 OR2_2033(g33065,g32008,g22068);
  OR2 OR2_2034(g34442,g34380,g18542);
  OR2 OR2_2035(g28513,g27276,g26123);
  OR2 OR2_2036(g31875,g31066,g21730);
  OR2 OR2_2037(g29643,g28192,g27145);
  OR2 OR2_2038(g34615,g34516,g18576);
  OR3 OR3_52(g33219,g32335,I30760,I30761);
  OR2 OR2_2039(g24262,g23387,g18315);
  OR2 OR2_2040(g28404,g27215,g15874);
  OR2 OR2_2041(g34720,g34694,g18134);
  OR2 OR2_2042(g34041,g33829,g18739);
  OR2 OR2_2043(g28717,g27482,g16701);
  OR2 OR2_2044(g30430,g29859,g21814);
  OR2 OR2_2045(g30493,g30198,g21989);
  OR2 OR2_2046(g28212,g27030,g27035);
  OR2 OR2_2047(g29260,g28315,g18604);
  OR2 OR2_2048(g25835,g25367,g23855);
  OR2 OR2_2049(g30465,g30164,g21936);
  OR2 OR2_2050(g34465,g34295,g18712);
  OR2 OR2_2051(g25586,g21678,g24156);
  OR2 OR2_2052(g34237,g32715,g33955);
  OR2 OR2_2053(g30340,g29377,g18245);
  OR2 OR2_2054(g29489,g28550,g27601);
  OR2 OR2_2055(g34035,g33721,g18714);
  OR2 OR2_2056(g29488,g28547,g27600);
  OR2 OR2_2057(g34806,g34763,g18595);
  OR2 OR2_2058(g23183,g19545,g15911);
  OR2 OR2_2059(g28723,g27490,g16706);
  OR2 OR2_2060(g33617,g33263,g24326);
  OR2 OR2_2061(g31915,g31520,g22001);
  OR2 OR2_2062(g25615,g24803,g18162);
  OR2 OR2_2063(g30517,g30244,g22038);
  OR2 OR2_2064(g28387,g27203,g15858);
  OR2 OR2_2065(g31277,g29570,g28285);
  OR2 OR2_2066(g25720,g25042,g18765);
  OR2 OR2_2067(g24247,g22623,g18259);
  OR2 OR2_2068(g33277,g32129,g29568);
  OR3 OR3_53(g14182,g11741,g11721,g753);
  OR2 OR2_2069(g15935,g13029,g10665);
  OR2 OR2_2070(g28097,g27682,g22005);
  OR2 OR2_2071(g28104,g27697,g22108);
  OR2 OR2_2072(g25746,g25217,g22063);
  OR2 OR2_2073(g28646,g27388,g16595);
  OR2 OR2_2074(g33595,g33368,g18489);
  OR2 OR2_2075(g32235,g31151,g29662);
  OR2 OR2_2076(g27562,g26102,g24703);
  OR2 OR2_2077(g33623,g33370,g18792);
  OR4 OR4_83(I30756,g32088,g32163,g32098,g32105);
  OR2 OR2_2078(g33037,g32177,g24310);
  OR2 OR2_2079(g30362,g30120,g18392);
  OR2 OR2_2080(g34193,g33809,g33814);
  OR2 OR2_2081(g24251,g22637,g18296);
  OR2 OR2_2082(g24272,g23056,g18629);
  OR2 OR2_2083(g31782,g30060,g30070);
  OR2 OR2_2084(g27290,g25926,g25928);
  OR2 OR2_2085(g28369,g27160,g25938);
  OR2 OR2_2086(g30523,g30245,g22069);
  OR2 OR2_2087(g33984,g33881,g18374);
  OR2 OR2_2088(g25684,g24983,g18643);
  OR2 OR2_2089(g29255,g28714,g18516);
  OR2 OR2_2090(g28368,g27158,g27184);
  OR2 OR2_2091(g26703,g24447,g10705);
  OR2 OR2_2092(g29270,g28258,g18635);
  OR2 OR2_2093(g32991,g32322,g18349);
  OR2 OR2_2094(g30475,g30220,g21946);
  OR2 OR2_2095(g34006,g33897,g18462);
  OR2 OR2_2096(g28850,g27557,g16869);
  OR2 OR2_2097(g33266,g32114,g29532);
  OR2 OR2_2098(g23574,g20093,g20108);
  OR2 OR2_2099(g13972,g11232,g11203);
  OR2 OR2_2100(g34727,g34655,g18213);
  OR2 OR2_2101(g26781,g24913,g24921);
  OR2 OR2_2102(g30437,g29876,g21846);
  OR2 OR2_2103(g26952,g26360,g24290);
  OR2 OR2_2104(g29294,g28645,g18779);
  OR2 OR2_2105(g29267,g28257,g18622);
  OR2 OR2_2106(g19619,g15712,g13080);
  OR2 OR2_2107(g8863,g1644,g1664);
  OR2 OR2_2108(g19557,g17123,g14190);
  OR3 OR3_54(I22830,g21429,g21338,g21307);
  OR2 OR2_2109(g27403,g25962,g24581);
  OR2 OR2_2110(g33589,g33340,g18469);
  OR2 OR2_2111(g30347,g29383,g18304);
  OR2 OR2_2112(g28716,g27481,g13887);
  OR2 OR2_2113(g34347,g25986,g34102);
  OR2 OR2_2114(g33588,g33334,g18468);
  OR2 OR2_2115(g34253,g34171,g24300);
  OR2 OR2_2116(g27226,g25872,g24436);
  OR2 OR2_2117(g28582,g27330,g26277);
  OR2 OR2_2118(g34600,g34538,g18182);
  OR2 OR2_2119(g24447,g10948,g22450);
  OR2 OR2_2120(g14387,g9086,g11048);
  OR2 OR2_2121(g34781,g33431,g34715);
  OR2 OR2_2122(g27551,g26091,g24675);
  OR2 OR2_2123(g27572,g26129,g24724);
  OR2 OR2_2124(g33119,g32420,g32428);
  OR2 OR2_2125(g28310,g27107,g15797);
  OR2 OR2_2126(g34236,g32650,g33954);
  OR2 OR2_2127(g30351,g30084,g18339);
  OR2 OR2_2128(g30372,g30110,g18446);
  OR2 OR2_2129(g25727,g25163,g22010);
  OR2 OR2_2130(g33118,g32413,g32418);
  OR2 OR2_2131(g34372,g26287,g34137);
  OR2 OR2_2132(g31864,g31271,g21703);
  OR2 OR2_2133(g33022,g32306,g21750);
  OR2 OR2_2134(g26422,g24774,g23104);
  OR2 OR2_2135(g31749,g29974,g29988);
  OR2 OR2_2136(g16052,g13060,g10724);
  OR2 OR2_2137(g7450,g1277,g1283);
  OR2 OR2_2138(g28050,g27692,g18165);
  OR2 OR2_2139(g33616,g33237,g24314);
  OR2 OR2_2140(g33313,g29649,g32171);
  OR2 OR2_2141(g30516,g30233,g22037);
  OR2 OR2_2142(g34264,g34081,g18701);
  OR2 OR2_2143(g28386,g27202,g13277);
  OR2 OR2_2144(g34790,g34774,g18151);
  OR2 OR2_2145(g31276,g29567,g28282);
  OR2 OR2_2146(g25703,g25087,g21922);
  OR2 OR2_2147(g28603,g27340,g26300);
  OR2 OR2_2148(g24246,g23372,g18257);
  OR2 OR2_2149(g33276,g32128,g29566);
  OR2 OR2_2150(g28096,g27988,g21997);
  OR2 OR2_2151(g32399,g31527,g30062);
  OR2 OR2_2152(g33053,g31967,g21974);
  OR2 OR2_2153(g31254,g25981,g29534);
  OR2 OR2_2154(g27980,g26105,g26131);
  OR2 OR2_2155(g33254,g32104,g29512);
  OR2 OR2_2156(g31900,g31484,g21908);
  OR2 OR2_2157(g31466,g26160,g29650);
  OR2 OR2_2158(g32398,g31526,g30061);
  OR3 OR3_55(I22267,g20236,g20133,g20111);
  OR2 OR2_2159(g25600,g24650,g18111);
  OR2 OR2_2160(g26913,g25848,g18225);
  OR2 OR2_2161(g28681,g27428,g16634);
  OR2 OR2_2162(g23405,g19791,g16245);
  OR2 OR2_2163(g29277,g28440,g18710);
  OR2 OR2_2164(g30422,g29795,g21806);
  OR2 OR2_2165(g33036,g32168,g24309);
  OR2 OR2_2166(g28429,g27228,g15913);
  OR2 OR2_2167(g33560,g33404,g18369);
  OR2 OR2_2168(g24355,g23799,g18824);
  OR2 OR2_2169(g28730,g27503,g13912);
  OR2 OR2_2170(g26905,g26397,g24222);
  OR4 OR4_84(g25821,g25482,g25456,g25417,g25377);
  OR2 OR2_2171(g28428,g27227,g15912);
  OR2 OR2_2172(g30542,g29337,g22088);
  OR2 OR2_2173(g30453,g29902,g21862);
  OR2 OR2_2174(g33064,g31993,g22067);
  OR2 OR2_2175(g19363,g17810,g14913);
  OR2 OR2_2176(g28690,g27436,g16641);
  OR2 OR2_2177(g34021,g33652,g18519);
  OR2 OR2_2178(g34453,g34410,g18666);
  OR2 OR2_2179(g27426,g25967,g24588);
  OR2 OR2_2180(g28549,g27304,g26233);
  OR2 OR2_2181(g24151,g18088,g21661);
  OR2 OR2_2182(g33733,g33105,g32012);
  OR2 OR2_2183(g32361,g29869,g31300);
  OR2 OR2_2184(g34726,g34665,g18212);
  OR2 OR2_2185(g28548,g27303,g26232);
  OR2 OR2_2186(g31874,g31016,g21729);
  OR2 OR2_2187(g30436,g29860,g21845);
  OR2 OR2_2188(g19486,g15589,g12979);
  OR2 OR2_2189(g34614,g34518,g18568);
  OR2 OR2_2190(g29266,g28330,g18621);
  OR2 OR2_2191(g34607,g34567,g15081);
  OR2 OR2_2192(g30530,g30224,g22076);
  OR2 OR2_2193(g28317,g27114,g15805);
  OR2 OR2_2194(g33009,g32273,g18458);
  OR2 OR2_2195(g34274,g27822,g34205);
  OR2 OR2_2196(g30346,g29381,g18303);
  OR2 OR2_2197(g25834,g25366,g23854);
  OR2 OR2_2198(g27024,g26826,g17692);
  OR4 OR4_85(I31849,g33483,g33484,g33485,g33486);
  OR2 OR2_2199(g33008,g32261,g18457);
  OR2 OR2_2200(g30464,g30152,g21935);
  OR2 OR2_2201(g32221,g31140,g29634);
  OR2 OR2_2202(g34464,g34340,g18687);
  OR2 OR2_2203(g31892,g31019,g21825);
  OR4 OR4_86(I31848,g33479,g33480,g33481,g33482);
  OR2 OR2_2204(g28057,g27033,g18218);
  OR2 OR2_2205(g34034,g33719,g18713);
  OR2 OR2_2206(g33555,g33355,g18357);
  OR2 OR2_2207(g34641,g34479,g18724);
  OR2 OR2_2208(g34797,g34747,g18574);
  OR2 OR2_2209(g25726,g25148,g22009);
  OR2 OR2_2210(g33570,g33420,g18405);
  OR2 OR2_2211(g31914,g31499,g22000);
  OR2 OR2_2212(g34292,g26853,g34223);
  OR2 OR2_2213(g28323,g27118,g15810);
  OR2 OR2_2214(g33914,g33305,g33311);
  OR2 OR2_2215(g34153,g33899,g33451);
  OR2 OR2_2216(g27126,g24378,g25787);
  OR2 OR2_2217(g25614,g24797,g18161);
  OR2 OR2_2218(g28533,g27291,g26203);
  OR2 OR2_2219(g31907,g31492,g21954);
  OR2 OR2_2220(g30409,g29842,g21768);
  OR2 OR2_2221(g27250,g25901,g15738);
  OR2 OR2_2222(g26891,g26652,g24197);
  OR2 OR2_2223(g24203,g22982,g18107);
  OR2 OR2_2224(g25607,g24773,g18118);
  OR2 OR2_2225(g10802,g7533,g1296);
  OR4 OR4_87(g15732,g13411,g13384,g13349,g11016);
  OR2 OR2_2226(g28775,g27537,g16806);
  OR2 OR2_2227(g30408,g29806,g21767);
  OR2 OR2_2228(g29864,g28272,g26086);
  OR2 OR2_2229(g34635,g34485,g18692);
  OR2 OR2_2230(g25593,g24716,g21707);
  OR2 OR2_2231(g33567,g33081,g18394);
  OR2 OR2_2232(g33594,g33421,g18485);
  OR2 OR2_2233(g32371,g29883,g31313);
  OR2 OR2_2234(g29313,g28284,g27270);
  OR2 OR2_2235(g24281,g23397,g18656);
  OR2 OR2_2236(g33238,g32048,g32051);
  OR2 OR2_2237(g26327,g8462,g24591);
  OR2 OR2_2238(g22225,g21332,g17654);
  OR2 OR2_2239(g29748,g28210,g28214);
  OR2 OR2_2240(g22708,g19266,g15711);
  OR2 OR2_2241(g29276,g28616,g18709);
  OR2 OR2_2242(g29285,g28639,g18750);
  OR2 OR2_2243(g29305,g28602,g18811);
  OR2 OR2_2244(g29254,g28725,g18512);
  OR3 OR3_56(g33176,g32198,I30734,I30735);
  OR2 OR2_2245(g16882,g13508,g11114);
  OR2 OR2_2246(g30474,g30208,g21945);
  OR2 OR2_2247(g25635,g24504,g18293);
  OR2 OR2_2248(g31883,g31132,g21777);
  OR2 OR2_2249(g30537,g30246,g22083);
  OR2 OR2_2250(g19587,g15700,g13046);
  OR4 OR4_88(I30331,g31672,g31710,g31021,g30937);
  OR2 OR2_2251(g34537,g34324,g34084);
  OR2 OR2_2252(g13794,g7396,g10684);
  OR2 OR2_2253(g34283,g26839,g34215);
  OR2 OR2_2254(g30492,g30188,g21988);
  OR2 OR2_2255(g34606,g34564,g15080);
  OR2 OR2_2256(g34303,g25768,g34045);
  OR2 OR2_2257(g28316,g27113,g15804);
  OR2 OR2_2258(g27581,g26161,g24750);
  OR2 OR2_2259(g27450,g2917,g26483);
  OR4 OR4_89(I30717,g31787,g32200,g31940,g31949);
  OR2 OR2_2260(g33577,g33405,g18430);
  OR2 OR2_2261(g30381,g30126,g18497);
  OR2 OR2_2262(g25575,g24139,g24140);
  OR2 OR2_2263(g28056,g27230,g18210);
  OR2 OR2_2264(g32359,g29867,g31298);
  OR2 OR2_2265(g27257,g25904,g24498);
  OR2 OR2_2266(g29166,g27653,g17153);
  OR2 OR2_2267(g25711,g25105,g21962);
  OR2 OR2_2268(g28611,g27348,g16485);
  OR2 OR2_2269(g24715,g22189,g22207);
  OR2 OR2_2270(g32358,g29866,g31297);
  OR2 OR2_2271(g34796,g34745,g18573);
  OR2 OR2_2272(g29892,g28300,g26120);
  OR2 OR2_2273(g27590,g26179,g24764);
  OR2 OR2_2274(g29476,g28108,g28112);
  OR2 OR2_2275(g29485,g28535,g27594);
  OR2 OR2_2276(g31906,g31477,g21953);
  OR2 OR2_2277(g30390,g29985,g18555);
  OR2 OR2_2278(g32344,g29804,g31266);
  OR2 OR2_2279(g31284,g29575,g28290);
  OR2 OR2_2280(g25606,g24761,g18117);
  OR2 OR2_2281(g28342,g27134,g15819);
  OR2 OR2_2282(g31304,g29594,g29608);
  OR3 OR3_57(g29914,g22531,g22585,I28147);
  OR2 OR2_2283(g21897,g20095,g15111);
  OR2 OR2_2284(g33622,g33366,g18791);
  OR2 OR2_2285(g33566,g33356,g18390);
  OR2 OR2_2286(g25750,g25543,g18802);
  OR2 OR2_2287(g26949,g26356,g24287);
  OR2 OR2_2288(g28650,g27391,g16598);
  OR2 OR2_2289(g30522,g29332,g22064);
  OR2 OR2_2290(g27150,g25804,g24400);
  OR2 OR2_2291(g34663,g32028,g34500);
  OR2 OR2_2292(g29239,g28427,g18297);
  OR2 OR2_2293(g26948,g26399,g24286);
  OR2 OR2_2294(g24354,g23775,g18823);
  OR2 OR2_2295(g27019,g26822,g14610);
  OR2 OR2_2296(g26904,g26393,g24221);
  OR2 OR2_2297(g29238,g28178,g18292);
  OR2 OR2_2298(g30483,g30241,g21979);
  OR2 OR2_2299(g30553,g30205,g22124);
  OR2 OR2_2300(g22901,g19384,g15745);
  OR2 OR2_2301(g28132,g27932,g27957);
  OR2 OR2_2302(g13997,g11029,g11036);
  OR2 OR2_2303(g29176,g27661,g17177);
  OR2 OR2_2304(g30536,g30234,g22082);
  OR2 OR2_2305(g26673,g24433,g10674);
  OR2 OR2_2306(g34040,g33818,g18737);
  OR2 OR2_2307(g33963,g33830,g18124);
  OR2 OR2_2308(g25663,g24666,g21788);
  OR2 OR2_2309(g34252,g34146,g18180);
  OR2 OR2_2310(g34621,g34517,g18583);
  OR2 OR2_2311(g28708,g27462,g16674);
  OR2 OR2_2312(g26933,g26808,g18551);
  OR2 OR2_2313(g28087,g27255,g18720);
  OR2 OR2_2314(g33576,g33401,g18423);
  OR2 OR2_2315(g33585,g33411,g18456);
  OR2 OR2_2316(g24211,g23572,g18138);
  OR2 OR2_2317(g28043,g27323,g21714);
  OR2 OR2_2318(g33554,g33407,g18353);
  OR2 OR2_2319(g32240,g24757,g31182);
  OR2 OR2_2320(g30397,g29747,g21756);
  OR4 OR4_90(I26742,g23430,g23445,g23458,g23481);
  OR2 OR2_2321(g33609,g33239,g18615);
  OR2 OR2_2322(g29501,g28583,g27634);
  OR2 OR2_2323(g33312,g29646,g32170);
  OR2 OR2_2324(g30509,g30210,g22030);
  OR2 OR2_2325(g33608,g33322,g18537);
  OR2 OR2_2326(g28069,g27564,g21865);
  OR2 OR2_2327(g33115,g32397,g32401);
  OR2 OR2_2328(g25702,g25068,g21921);
  OR2 OR2_2329(g25757,g25132,g22104);
  OR2 OR2_2330(g28774,g27536,g16804);
  OR2 OR2_2331(g30508,g30199,g22029);
  OR2 OR2_2332(g31921,g31508,g22046);
  OR2 OR2_2333(g28068,g27310,g21838);
  OR2 OR2_2334(g32981,g32425,g18206);
  OR2 OR2_2335(g28375,g27183,g15851);
  OR2 OR2_2336(g33052,g31961,g21973);
  OR2 OR2_2337(g34634,g34483,g18691);
  OR2 OR2_2338(g25621,g24523,g18205);
  OR2 OR2_2339(g31745,g29959,g29973);
  OR2 OR2_2340(g21896,g20084,g15110);
  OR2 OR2_2341(g24250,g22633,g18295);
  OR2 OR2_2342(g26912,g25946,g18209);
  OR2 OR2_2343(g27231,g25873,g15699);
  OR2 OR2_2344(g29284,g28554,g18747);
  OR2 OR2_2345(g32395,g31523,g30049);
  OR2 OR2_2346(g24339,g23690,g18756);
  OR2 OR2_2347(g33973,g33840,g18344);
  OR2 OR2_2348(g29304,g28588,g18810);
  OR2 OR2_2349(g32262,g31186,g29710);
  OR2 OR2_2350(g23716,g9194,g20905);
  OR2 OR2_2351(g25673,g24727,g21830);
  OR2 OR2_2352(g32990,g32281,g18341);
  OR3 OR3_58(I18417,g14444,g14414,g14392);
  OR2 OR2_2353(g24338,g23658,g18755);
  OR2 OR2_2354(g11370,g8807,g550);
  OR2 OR2_2355(g30452,g29891,g21861);
  OR2 OR2_2356(g34452,g34401,g18665);
  OR2 OR2_2357(g13858,g209,g10685);
  OR2 OR2_2358(g33732,g33104,g32011);
  OR2 OR2_2359(g30311,g28265,g27265);
  OR3 OR3_59(g24968,g22360,g22409,g23389);
  OR2 OR2_2360(g25634,g24559,g18284);
  OR2 OR2_2361(g31761,g30009,g30028);
  OR2 OR2_2362(g33692,g32400,g33428);
  OR2 OR2_2363(g19475,g16930,g14126);
  OR2 OR2_2364(g27456,g25978,g24607);
  OR2 OR2_2365(g26396,g24762,g23062);
  OR2 OR2_2366(g28545,g27301,g26230);
  OR2 OR2_2367(g28078,g27140,g21880);
  OR2 OR2_2368(g33013,g32283,g18484);
  OR2 OR2_2369(g22669,g7763,g19525);
  OR2 OR2_2370(g32247,g31168,g29686);
  OR3 OR3_60(I18543,g14568,g14540,g14516);
  OR2 OR2_2371(g28086,g27268,g18702);
  OR2 OR2_2372(g32389,g31496,g29966);
  OR2 OR2_2373(g30350,g30118,g18334);
  OR2 OR2_2374(g34350,g26048,g34106);
  OR2 OR2_2375(g33539,g33245,g18178);
  OR2 OR2_2376(g32388,g31495,g29962);
  OR2 OR2_2377(g33005,g32260,g18432);
  OR2 OR2_2378(g27596,g26207,g24775);
  OR2 OR2_2379(g11025,g2980,g7831);
  OR2 OR2_2380(g28817,g27548,g16845);
  OR2 OR2_2381(g33538,g33252,g18144);
  OR2 OR2_2382(g28322,g27117,g15809);
  OR2 OR2_2383(g27243,g25884,g24475);
  OR2 OR2_2384(g30396,g29856,g21755);
  OR2 OR2_2385(g32251,g30599,g29352);
  OR2 OR2_2386(g13540,g10822,g10827);
  OR2 OR2_2387(g27431,g24582,g25977);
  OR2 OR2_2388(g20202,g16211,g13507);
  OR2 OR2_2389(g34731,g34662,g18272);
  OR2 OR2_2390(g29484,g28124,g22191);
  OR2 OR2_2391(g24202,g22899,g18106);
  OR2 OR2_2392(g26929,g26635,g18543);
  OR2 OR2_2393(g24257,g22938,g18310);
  OR2 OR2_2394(g30413,g30001,g21772);
  OR2 OR2_2395(g24496,g24008,g21557);
  OR2 OR2_2396(g31241,g25959,g29510);
  OR2 OR2_2397(g26928,g26713,g18541);
  OR4 OR4_91(g17488,g14361,g14335,g11954,I18417);
  OR2 OR2_2398(g25592,g24672,g21706);
  OR2 OR2_2399(g25756,g25112,g22103);
  OR2 OR2_2400(g28561,g27312,g26250);
  OR2 OR2_2401(g28295,g27094,g15783);
  OR2 OR2_2402(g28680,g27427,g16633);
  OR2 OR2_2403(g32997,g32269,g18378);
  OR2 OR2_2404(g30405,g29767,g21764);
  OR2 OR2_2405(g16173,g8796,g13464);
  OR2 OR2_2406(g34405,g34183,g25103);
  OR2 OR2_2407(g33235,g32040,g30982);
  OR2 OR2_2408(g23317,g19715,g16191);
  OR3 OR3_61(I22852,g21459,g21350,g21339);
  OR2 OR2_2409(g29813,g26020,g28261);
  OR2 OR2_2410(g22679,g19145,g15701);
  OR2 OR2_2411(g23129,g19500,g15863);
  OR2 OR2_2412(g13699,g10921,g10947);
  OR2 OR2_2413(g34020,g33904,g18514);
  OR2 OR2_2414(g25731,g25128,g22014);
  OR2 OR2_2415(g28631,g27372,g16534);
  OR4 OR4_92(I28567,g29204,g29205,g29206,g29207);
  OR3 OR3_62(I24117,g23088,g23154,g23172);
  OR2 OR2_2416(g32360,g29868,g31299);
  OR2 OR2_2417(g16506,g13294,g10966);
  OR2 OR2_2418(g15789,g10819,g13211);
  OR4 OR4_93(I30261,g29385,g31376,g30735,g30825);
  OR2 OR2_2419(g34046,g33906,g33908);
  OR2 OR2_2420(g31882,g31115,g21776);
  OR2 OR2_2421(g33991,g33885,g18400);
  OR2 OR2_2422(g14078,g10776,g8703);
  OR2 OR2_2423(g20196,g16207,g13497);
  OR2 OR2_2424(g25691,g24536,g21890);
  OR2 OR2_2425(g27487,g25990,g24629);
  OR2 OR2_2426(g34282,g26838,g34214);
  OR2 OR2_2427(g23298,g19693,g16179);
  OR2 OR2_2428(g30357,g30107,g18366);
  OR2 OR2_2429(g28309,g27106,g15796);
  OR2 OR2_2430(g32220,g31139,g29633);
  OR2 OR2_2431(g26881,g26629,g24187);
  OR2 OR2_2432(g16927,g13524,g11126);
  OR2 OR2_2433(g25929,g24395,g22193);
  OR2 OR2_2434(g28308,g27105,g15795);
  OR2 OR2_2435(g27278,g15786,g25921);
  OR2 OR2_2436(g29692,g28197,g10873);
  OR2 OR2_2437(g24457,g10902,g22400);
  OR2 OR2_2438(g14977,g10776,g8703);
  OR2 OR2_2439(g25583,g21666,g24153);
  OR2 OR2_2440(g33584,g33406,g18449);
  OR2 OR2_2441(g34640,g34487,g18723);
  OR2 OR2_2442(g19274,g17753,g14791);
  OR2 OR2_2443(g19593,g17145,g14210);
  OR2 OR2_2444(g34803,g34758,g18590);
  OR2 OR2_2445(g28816,g27547,g16843);
  OR2 OR2_2446(g20077,g16025,g13320);
  OR2 OR2_2447(g23261,g19660,g16125);
  OR2 OR2_2448(g26890,g26630,g24196);
  OR2 OR2_2449(g28687,g27434,g16638);
  OR2 OR2_2450(g29539,g2864,g28220);
  OR2 OR2_2451(g32355,g29855,g31286);
  OR2 OR2_2452(g34881,g34866,g18187);
  OR2 OR2_2453(g24256,g22873,g18309);
  OR2 OR2_2454(g32370,g29882,g31312);
  OR2 OR2_2455(g28374,g27181,g15850);
  OR2 OR2_2456(g24280,g23292,g15109);
  OR2 OR2_2457(g25743,g25110,g22058);
  OR2 OR2_2458(g28643,g27386,g16592);
  OR2 OR2_2459(g27937,g14506,g26793);
  OR2 OR2_2460(g32996,g32256,g18377);
  OR2 OR2_2461(g34027,g33718,g18683);
  OR2 OR2_2462(g29241,g28638,g18332);
  OR2 OR2_2463(g13385,g11967,g9479);
  ND2 NAND2_0(g11980,I14817,I14818);
  ND2 NAND2_1(g13889,g11566,g11435);
  ND2 NAND2_2(g13980,g10295,g11435);
  ND2 NAND2_3(g12169,g9804,g5448);
  ND2 NAND2_4(I22761,g11939,I22760);
  ND2 NAND2_5(I13443,g262,I13442);
  ND2 NAND2_6(I14185,g8442,g3470);
  ND4 NAND4_0(g16719,g3243,g13700,g3310,g11350);
  ND2 NAND2_7(I14518,g661,I14516);
  ND4 NAND4_1(g10224,g6661,g6704,g6675,g6697);
  ND2 NAND2_8(g17595,g8616,g14367);
  ND2 NAND2_9(g22984,g20114,g2868);
  ND2 NAND2_10(I12346,g3111,I12344);
  ND2 NAND2_11(g12478,I15299,I15300);
  ND4 NAND4_2(g21432,g17790,g14820,g17761,g14780);
  ND3 NAND3_0(g28830,g27886,g7451,g7369);
  ND2 NAND2_12(I14883,g9500,g5489);
  ND2 NAND2_13(g19474,g11609,g17794);
  ND2 NAND2_14(g11426,g8742,g4878);
  ND2 NAND2_15(g11190,g8539,g3447);
  ND2 NAND2_16(g9852,g3684,g4871);
  ND2 NAND2_17(g23342,g6928,g21163);
  ND2 NAND2_18(g27223,I25908,I25909);
  ND2 NAND2_19(I15089,g2393,I15087);
  ND2 NAND2_20(g22853,g20219,g2922);
  ND2 NAND2_21(g25003,g21353,g23462);
  ND2 NAND2_22(I15088,g9832,I15087);
  ND2 NAND2_23(g24916,g19450,g23154);
  ND2 NAND2_24(g25779,g19694,g24362);
  ND2 NAND2_25(g12084,g2342,g8211);
  ND3 NAND3_1(g28270,g10504,g26105,g26987);
  ND2 NAND2_26(g22836,g18918,g2852);
  ND2 NAND2_27(g21330,g11401,g17157);
  ND2 NAND2_28(g20076,g13795,g16521);
  ND4 NAND4_3(g21365,g15744,g13119,g15730,g13100);
  ND2 NAND2_29(g23132,g8155,g19932);
  ND2 NAND2_30(I22683,g11893,g21434);
  ND2 NAND2_31(g28938,g27796,g8205);
  ND2 NAND2_32(g9825,I13391,I13392);
  ND2 NAND2_33(g7201,I11865,I11866);
  ND4 NAND4_4(g15719,g5256,g14490,g5335,g9780);
  ND3 NAND3_2(g27654,g164,g26598,g23042);
  ND2 NAND2_34(g22864,g7780,g21156);
  ND2 NAND2_35(I20165,g16246,g990);
  ND2 NAND2_36(g14489,g12126,g5084);
  ND2 NAND2_37(g29082,g27837,g9694);
  ND2 NAND2_38(g25233,g20838,g23623);
  ND2 NAND2_39(g24942,g20039,g23172);
  ND2 NAND2_40(I26459,g26576,g14306);
  ND3 NAND3_3(g15832,g7903,g7479,g13256);
  ND4 NAND4_5(g14830,g6605,g12211,g6723,g12721);
  ND2 NAND2_41(I32431,g34056,g34051);
  ND2 NAND2_42(g9972,I13510,I13511);
  ND2 NAND2_43(I20222,g16272,I20221);
  ND3 NAND3_4(g17748,g562,g14708,g12323);
  ND2 NAND2_44(g11969,g7252,g1636);
  ND2 NAND2_45(g20734,g14408,g17312);
  ND3 NAND3_5(g28837,g27800,g7374,g2197);
  ND2 NAND2_46(I25244,g24744,I25242);
  ND3 NAND3_6(g11968,g837,g9334,g9086);
  ND4 NAND4_6(g13968,g3913,g11255,g4031,g11631);
  ND2 NAND2_47(g15045,g12716,g7142);
  ND2 NAND2_48(g12423,I15242,I15243);
  ND4 NAND4_7(g27587,g24917,g25018,g24918,g26857);
  ND2 NAND2_49(g20838,g5041,g17284);
  ND2 NAND2_50(g13855,g4944,g11804);
  ND3 NAND3_7(g19483,g15969,g10841,g10922);
  ND2 NAND2_51(g10610,g7462,g7490);
  ND2 NAND2_52(g11411,g9713,g3625);
  ND2 NAND2_53(I13110,g5808,I13109);
  ND2 NAND2_54(g22642,g7870,g19560);
  ND2 NAND2_55(g12587,g7497,g6315);
  ND2 NAND2_56(g13870,g11773,g4732);
  ND4 NAND4_8(g13527,g182,g168,g203,g12812);
  ND2 NAND2_57(g23810,I22973,I22974);
  ND2 NAND2_58(g20619,g14317,g17217);
  ND4 NAND4_9(g16628,g3602,g11207,g3618,g13902);
  ND2 NAND2_59(I23119,g20076,I23118);
  ND4 NAND4_10(g10124,g5276,g5320,g5290,g5313);
  ND2 NAND2_60(g12000,g8418,g2610);
  ND2 NAND2_61(I23118,g20076,g417);
  ND2 NAND2_62(g22874,g18918,g2844);
  ND2 NAND2_63(g10939,g7352,g1459);
  ND2 NAND2_64(g13867,g11312,g8449);
  ND4 NAND4_11(g14686,g5268,g12059,g5276,g12239);
  ND2 NAND2_65(I12840,g4222,g4235);
  ND2 NAND2_66(g29049,g9640,g27779);
  ND4 NAND4_12(g16776,g3945,g13772,g4012,g11419);
  ND2 NAND2_67(g13315,g1459,g10715);
  ND2 NAND2_68(g11707,g8718,g4864);
  ND2 NAND2_69(I18530,g1811,I18529);
  ND2 NAND2_70(g20039,g11250,g17794);
  ND2 NAND2_71(I14609,g8993,g8678);
  ND2 NAND2_72(I13334,g1687,g1691);
  ND2 NAND2_73(g13257,g1389,g10544);
  ND2 NAND2_74(g29004,g27933,g8330);
  ND4 NAND4_13(g21459,g17814,g14854,g17605,g17581);
  ND2 NAND2_75(g11979,g9861,g5452);
  ND3 NAND3_8(g13496,g1351,g11336,g11815);
  ND3 NAND3_9(g11590,g6928,g3990,g4049);
  ND3 NAND3_10(g12639,g10194,g6682,g6732);
  ND2 NAND2_76(g22712,g18957,g2864);
  ND2 NAND2_77(g23010,g20516,g2984);
  ND2 NAND2_78(g7897,I12288,I12289);
  ND2 NAND2_79(g24601,g22957,g2965);
  ND2 NAND2_80(g13986,g10323,g11747);
  ND2 NAND2_81(g12293,g7436,g5283);
  ND2 NAND2_82(g24677,g22957,g2975);
  ND2 NAND2_83(g12638,g7514,g6661);
  ND2 NAND2_84(g24975,g21388,g23363);
  ND4 NAND4_14(g10160,g5623,g5666,g5637,g5659);
  ND4 NAND4_15(g17712,g5599,g14425,g5666,g12301);
  ND3 NAND3_11(g12416,g10133,g7064,g10166);
  ND2 NAND2_85(g14160,g11626,g8958);
  ND3 NAND3_12(g28853,g27742,g1636,g7252);
  ND4 NAND4_16(g13067,g5240,g12059,g5331,g9780);
  ND2 NAND2_86(g28167,g925,g27046);
  ND2 NAND2_87(I18635,g14713,I18633);
  ND2 NAND2_88(g10617,g10151,g9909);
  ND3 NAND3_13(g16319,g8224,g8170,g13736);
  ND2 NAND2_89(I32187,g33661,I32185);
  ND2 NAND2_90(I12252,g1124,I12251);
  ND2 NAND2_91(g14915,g12553,g10266);
  ND2 NAND2_92(g22941,g20219,g2970);
  ND2 NAND2_93(I17406,g1472,I17404);
  ND2 NAND2_94(g12578,g7791,g10341);
  ND4 NAND4_17(g27586,g24924,g24916,g24905,g26863);
  ND2 NAND2_95(g12014,g7197,g703);
  ND2 NAND2_96(g14075,g11658,g11527);
  ND3 NAND3_14(g15591,g4332,g4322,g13202);
  ND3 NAND3_15(g28864,g27886,g7411,g1996);
  ND2 NAND2_97(g10623,g10181,g9976);
  ND4 NAND4_18(g17675,g5252,g14399,g5320,g12239);
  ND2 NAND2_98(g23656,I22800,I22801);
  ND2 NAND2_99(g21353,g11467,g17157);
  ND2 NAND2_100(I13751,g4584,I13749);
  ND2 NAND2_101(g14782,g12755,g10491);
  ND2 NAND2_102(I14400,g3654,I14398);
  ND2 NAND2_103(g12116,g2051,g8255);
  ND2 NAND2_104(g14984,g7812,g12680);
  ND4 NAND4_19(g13866,g3239,g11194,g3321,g11519);
  ND2 NAND2_105(I18537,g2236,I18536);
  ND3 NAND3_16(g16281,g4754,g13937,g12054);
  ND3 NAND3_17(g28900,g27886,g7451,g2040);
  ND2 NAND2_106(g14822,g12755,g12632);
  ND2 NAND2_107(g14170,g11715,g11537);
  ND3 NAND3_18(g15844,g14714,g9340,g12378);
  ND2 NAND2_108(I22972,g9657,g19638);
  ND4 NAND4_20(g21364,g15787,g15781,g15753,g13131);
  ND2 NAND2_109(I13391,g1821,I13390);
  ND3 NAND3_19(g13256,g11846,g11294,g11812);
  ND2 NAND2_110(I13510,g2089,I13509);
  ND2 NAND2_111(g11923,I14734,I14735);
  ND2 NAND2_112(g12340,g4888,g8984);
  ND2 NAND2_113(g12035,g10000,g6144);
  ND2 NAND2_114(g13923,g11692,g11527);
  ND2 NAND2_115(I15300,g1982,I15298);
  ND2 NAND2_116(g9830,I13402,I13403);
  ND2 NAND2_117(g20186,g16926,g8177);
  ND2 NAND2_118(g20676,g14379,g17287);
  ND2 NAND2_119(g21289,g14616,g17493);
  ND2 NAND2_120(I12205,g1135,I12203);
  ND2 NAND2_121(g13102,g7523,g10759);
  ND3 NAND3_20(g25429,g22417,g1917,g8302);
  ND2 NAND2_122(g23309,g6905,g21024);
  ND3 NAND3_21(g28874,g27907,g7424,g2421);
  ND2 NAND2_123(g29121,g9755,g27886);
  ND2 NAND2_124(g21288,g14616,g17492);
  ND2 NAND2_125(g7582,g1361,g1373);
  ND2 NAND2_126(I13442,g262,g239);
  ND3 NAND3_22(g13066,g4430,g7178,g10590);
  ND4 NAND4_21(g24936,g20186,g20173,g23379,g14029);
  ND3 NAND3_23(g31262,g767,g29916,g11679);
  ND2 NAND2_127(g10022,g6474,g6466);
  ND2 NAND2_128(g14864,g7791,g10421);
  ND2 NAND2_129(g8769,g691,g714);
  ND2 NAND2_130(g7227,g4584,g4593);
  ND2 NAND2_131(I32186,g33665,I32185);
  ND2 NAND2_132(g12523,g7563,g6346);
  ND3 NAND3_24(g28892,g27779,g1772,g7275);
  ND2 NAND2_133(g13854,g4765,g11797);
  ND2 NAND2_134(g11511,I14481,I14482);
  ND2 NAND2_135(I14991,g9685,g6527);
  ND2 NAND2_136(g8967,g4264,g4258);
  ND4 NAND4_22(g13511,g182,g174,g203,g12812);
  ND2 NAND2_137(g20216,I20487,I20488);
  ND3 NAND3_25(g14254,g11968,g11933,g11951);
  ND3 NAND3_26(g28914,g27937,g7462,g2555);
  ND2 NAND2_138(g29134,g9762,g27907);
  ND3 NAND3_27(g28907,g27858,g2361,g2287);
  ND2 NAND2_139(g12222,g8310,g2028);
  ND2 NAND2_140(g29028,g27933,g8381);
  ND2 NAND2_141(g22852,g18957,g2856);
  ND2 NAND2_142(g14101,g11653,g11729);
  ND2 NAND2_143(g25002,g19474,g23154);
  ND2 NAND2_144(I29297,g12117,I29295);
  ND3 NAND3_28(g14177,g11741,g11721,g753);
  ND2 NAND2_145(g11480,g10323,g8906);
  ND2 NAND2_146(I26460,g26576,I26459);
  ND2 NAND2_147(I22946,g19620,I22944);
  ND2 NAND2_148(I18536,g2236,g14642);
  ND2 NAND2_149(I15287,g10061,g6697);
  ND2 NAND2_150(I14206,g3821,I14204);
  ND4 NAND4_23(g16956,g3925,g13824,g4019,g11631);
  ND2 NAND2_151(I26093,g26055,g13539);
  ND2 NAND2_152(I15307,g10116,I15306);
  ND2 NAND2_153(g23195,g20136,g37);
  ND2 NAND2_154(g13307,g1116,g10695);
  ND2 NAND2_155(I15243,g6351,I15241);
  ND4 NAND4_24(g16181,g13475,g13495,g13057,g13459);
  ND2 NAND2_156(g12351,I15194,I15195);
  ND2 NAND2_157(g24814,g20011,g23167);
  ND2 NAND2_158(g22312,g907,g19063);
  ND3 NAND3_29(g28935,g27800,g2227,g7328);
  ND2 NAND2_159(g24807,I23979,I23980);
  ND2 NAND2_160(I15341,g10154,I15340);
  ND2 NAND2_161(g14665,g12604,g12798);
  ND2 NAND2_162(g24974,g21301,g23363);
  ND2 NAND2_163(g31997,g22306,g30580);
  ND2 NAND2_164(g14008,g11610,g11435);
  ND2 NAND2_165(I14399,g8542,I14398);
  ND2 NAND2_166(I22760,g11939,g21434);
  ND2 NAND2_167(g9258,I13044,I13045);
  ND2 NAND2_168(g22921,g20219,g2950);
  ND3 NAND3_30(g15715,g336,g305,g13385);
  ND2 NAND2_169(g17312,g7297,g14248);
  ND2 NAND2_170(g25995,g24621,g22853);
  ND2 NAND2_171(g14892,g12700,g12515);
  ND4 NAND4_25(g17608,g5953,g12067,g5969,g14701);
  ND2 NAND2_172(I14398,g8542,g3654);
  ND2 NAND2_173(g15572,g12969,g7219);
  ND2 NAND2_174(I18634,g2504,I18633);
  ND2 NAND2_175(I15335,g2116,I15333);
  ND2 NAND2_176(g34056,I31984,I31985);
  ND4 NAND4_26(g14570,g3933,g11255,g4023,g8595);
  ND2 NAND2_177(g11993,g1894,g8302);
  ND4 NAND4_27(g13993,g3961,g11255,g3969,g11419);
  ND2 NAND2_178(I23963,g13631,I23961);
  ND2 NAND2_179(g9975,I13519,I13520);
  ND2 NAND2_180(g21124,g5731,g17393);
  ND2 NAND2_181(I14332,g9966,I14330);
  ND2 NAND2_182(g13667,g3723,g11119);
  ND4 NAND4_28(g13131,g6243,g12101,g6377,g10003);
  ND2 NAND2_183(g10567,g1862,g7405);
  ND2 NAND2_184(g20007,g11512,g17794);
  ND2 NAND2_185(I23585,g22409,g4332);
  ND4 NAND4_29(g28349,g27074,g24770,g27187,g19644);
  ND2 NAND2_186(g29719,g28406,g13739);
  ND2 NAND2_187(g21294,g11324,g17157);
  ND3 NAND3_31(g25498,g22498,g2610,g8418);
  ND2 NAND2_188(g28906,g27796,g8150);
  ND2 NAND2_189(g13210,g7479,g10521);
  ND2 NAND2_190(g34650,I32757,I32758);
  ND4 NAND4_30(g16625,g3203,g13700,g3274,g11519);
  ND4 NAND4_31(g17732,g3937,g13824,g4012,g13933);
  ND4 NAND4_32(g10185,g5969,g6012,g5983,g6005);
  ND2 NAND2_191(g11443,g9916,g3649);
  ND2 NAND2_192(g12436,I15263,I15264);
  ND2 NAND2_193(g11279,g8504,g3443);
  ND4 NAND4_33(g14519,g3889,g11225,g4000,g8595);
  ND2 NAND2_194(I29296,g29495,I29295);
  ND2 NAND2_195(g14675,g12317,g9898);
  ND2 NAND2_196(I25219,g482,g24718);
  ND4 NAND4_34(g27593,g24972,g24950,g24906,g26861);
  ND2 NAND2_197(I26419,g14247,I26417);
  ND2 NAND2_198(I22755,g21434,I22753);
  ND2 NAND2_199(g12073,g10058,g6490);
  ND2 NAND2_200(g14154,g11669,g8958);
  ND4 NAND4_35(g17761,g6291,g14529,g6358,g12423);
  ND2 NAND2_201(I26418,g26519,I26417);
  ND2 NAND2_202(g13469,g4983,g10862);
  ND2 NAND2_203(g25432,g12374,g22384);
  ND2 NAND2_204(g10935,g1459,g7352);
  ND2 NAND2_205(g14637,g12255,g9815);
  ND2 NAND2_206(I15306,g10116,g2407);
  ND2 NAND2_207(g16296,g9360,g13501);
  ND2 NAND2_208(g25271,I24462,I24463);
  ND2 NAND2_209(g7133,I11825,I11826);
  ND3 NAND3_32(g12464,g10169,g7087,g10191);
  ND2 NAND2_210(g7846,g4843,g4878);
  ND4 NAND4_36(g12797,g10275,g7655,g7643,g7627);
  ND2 NAND2_211(I22794,g21434,I22792);
  ND2 NAND2_212(I22845,g12113,I22844);
  ND2 NAND2_213(g7803,I12204,I12205);
  ND2 NAND2_214(g31950,g7285,g30573);
  ND2 NAND2_215(g12292,g4698,g8933);
  ND2 NAND2_216(g9461,I13140,I13141);
  ND2 NAND2_217(g12153,g2610,g8330);
  ND2 NAND2_218(g25199,I24364,I24365);
  ND2 NAND2_219(I22899,g12193,g21228);
  ND2 NAND2_220(g8829,g5011,g4836);
  ND2 NAND2_221(g11975,g8267,g8316);
  ND2 NAND2_222(I12204,g1094,I12203);
  ND3 NAND3_33(g19513,g15969,g10841,g10922);
  ND2 NAND2_223(g23617,I22761,I22762);
  ND2 NAND2_224(g15024,g12780,g10421);
  ND2 NAND2_225(I20205,g11147,I20203);
  ND2 NAND2_226(g12136,I14992,I14993);
  ND2 NAND2_227(I22719,g21434,I22717);
  ND2 NAND2_228(g9904,I13443,I13444);
  ND4 NAND4_37(g13143,g10695,g7661,g979,g1061);
  ND2 NAND2_229(I13453,g1955,I13452);
  ND2 NAND2_230(I22718,g11916,I22717);
  ND3 NAND3_34(g33394,g10159,g4474,g32426);
  ND2 NAND2_231(g11169,I14229,I14230);
  ND2 NAND2_232(I29315,g12154,I29313);
  ND2 NAND2_233(I15168,g9823,I15166);
  ND2 NAND2_234(g13884,g11797,g4727);
  ND3 NAND3_35(g11410,g6875,g6895,g8696);
  ND2 NAND2_235(g23623,g9364,g20717);
  ND2 NAND2_236(g9391,I13110,I13111);
  ND2 NAND2_237(I15363,g10182,g2675);
  ND2 NAND2_238(g8124,I12402,I12403);
  ND2 NAND2_239(g24362,g21370,g22136);
  ND3 NAND3_36(g11479,g6875,g3288,g3347);
  ND2 NAND2_240(g23782,g2741,g21062);
  ND2 NAND2_241(g13666,g11190,g8441);
  ND4 NAND4_38(g13479,g12686,g12639,g12590,g12526);
  ND2 NAND2_242(g8069,I12373,I12374);
  ND2 NAND2_243(I32517,g34424,I32516);
  ND2 NAND2_244(g13217,g4082,g10808);
  ND2 NAND2_245(g10622,g10178,g9973);
  ND2 NAND2_246(g10566,g7315,g7356);
  ND4 NAND4_39(g13478,g12511,g12460,g12414,g12344);
  ND2 NAND2_247(I13565,g2648,I13564);
  ND2 NAND2_248(I13464,g2384,I13462);
  ND3 NAND3_37(g13486,g10862,g4983,g4966);
  ND2 NAND2_249(g25258,I24439,I24440);
  ND2 NAND2_250(g23266,g18918,g2894);
  ND4 NAND4_40(g13580,g11849,g7503,g7922,g10544);
  ND2 NAND2_251(g10653,g10204,g10042);
  ND2 NAND2_252(g14139,g11626,g11584);
  ND4 NAND4_41(g16741,g3207,g13765,g3303,g11519);
  ND2 NAND2_253(I14789,g9891,I14788);
  ND2 NAND2_254(g23167,g8219,g19981);
  ND4 NAND4_42(g13084,g5587,g12093,g5677,g9864);
  ND3 NAND3_38(g28973,g27907,g2465,g7387);
  ND4 NAND4_43(g14636,g5595,g12029,g5677,g12563);
  ND2 NAND2_255(I14788,g9891,g6167);
  ND4 NAND4_44(g14333,g12042,g12014,g11990,g11892);
  ND2 NAND2_256(I17462,g1300,I17460);
  ND4 NAND4_45(g21401,g17755,g14730,g17712,g14695);
  ND4 NAND4_46(g27796,g21228,g25263,g26424,g26171);
  ND4 NAND4_47(g20236,g16875,g14014,g16625,g16604);
  ND2 NAND2_257(g12796,g4467,g6961);
  ND2 NAND2_258(g9654,g2485,g2453);
  ND3 NAND3_39(g15867,g14714,g9417,g9340);
  ND3 NAND3_40(g25337,g22342,g1648,g8187);
  ND2 NAND2_259(g28934,g27882,g14641);
  ND4 NAND4_48(g14664,g5220,g12059,g5339,g12497);
  ND4 NAND4_49(g16196,g13496,g13513,g13079,g13476);
  ND4 NAND4_50(g11676,g358,g8944,g376,g385);
  ND3 NAND3_41(g34545,g11679,g794,g34354);
  ND2 NAND2_260(I22871,g12150,g21228);
  ND2 NAND2_261(g11953,g8195,g8241);
  ND2 NAND2_262(g13676,g11834,g11283);
  ND2 NAND2_263(g23616,I22754,I22755);
  ND2 NAND2_264(g29355,g24383,g28109);
  ND2 NAND2_265(g15581,g7232,g12999);
  ND2 NAND2_266(g10585,g1996,g7451);
  ND2 NAND2_267(g9595,g2351,g2319);
  ND2 NAND2_268(g23748,I22872,I22873);
  ND2 NAND2_269(I14291,g3835,I14289);
  ND2 NAND2_270(g11936,g8241,g1783);
  ND2 NAND2_271(I15334,g10152,I15333);
  ND2 NAND2_272(g12192,g8267,g2319);
  ND2 NAND2_273(g10609,g10111,g9826);
  ND2 NAND2_274(I13109,g5808,g5813);
  ND2 NAND2_275(g22940,g18918,g2860);
  ND2 NAND2_276(I12097,g1339,I12096);
  ND2 NAND2_277(g25425,g20081,g23172);
  ND3 NAND3_42(g12522,g10133,g5990,g6040);
  ND2 NAND2_278(g23809,I22966,I22967);
  ND4 NAND4_51(g17744,g6303,g14529,g6373,g12672);
  ND2 NAND2_279(I17447,g13336,I17446);
  ND3 NAND3_43(g28207,g12546,g26131,g27977);
  ND3 NAND3_44(g17399,g9626,g9574,g14535);
  ND2 NAND2_280(g14921,g12492,g10266);
  ND4 NAND4_52(g15741,g5244,g14490,g5320,g14631);
  ND2 NAND2_281(I32516,g34424,g34422);
  ND2 NAND2_282(g9629,g6462,g6466);
  ND2 NAND2_283(I13750,g4608,I13749);
  ND2 NAND2_284(g14813,g7766,g12824);
  ND2 NAND2_285(g11543,g9714,g3969);
  ND2 NAND2_286(I12850,g4277,I12848);
  ND4 NAND4_53(g13909,g11396,g8847,g11674,g8803);
  ND2 NAND2_287(g23733,g20751,g11178);
  ND4 NAND4_54(g15735,g5547,g14425,g5659,g9864);
  ND3 NAND3_45(g15877,g14833,g9340,g12543);
  ND2 NAND2_288(g9800,g5436,g5428);
  ND4 NAND4_55(g14674,g5941,g12067,g6023,g12614);
  ND3 NAND3_46(g11117,g8087,g8186,g8239);
  ND3 NAND3_47(g29025,g27937,g2629,g7462);
  ND2 NAND2_289(g13000,g7228,g10598);
  ND2 NAND2_290(I22754,g11937,I22753);
  ND2 NAND2_291(g29540,g28336,g13464);
  ND2 NAND2_292(g23630,g20739,g11123);
  ND3 NAND3_48(g22833,g1193,g19560,g10666);
  ND2 NAND2_293(g15695,g1266,g13125);
  ND2 NAND2_294(g25532,g21360,g23363);
  ND2 NAND2_295(g15018,g12739,g12515);
  ND2 NAND2_296(I13390,g1821,g1825);
  ND2 NAND2_297(g14732,g12662,g12515);
  ND2 NAND2_298(g24905,g534,g23088);
  ND2 NAND2_299(I15242,g10003,I15241);
  ND2 NAND2_300(g19857,g13628,g16296);
  ND2 NAND2_301(g17500,g14573,g14548);
  ND2 NAND2_302(I15123,g2102,I15121);
  ND2 NAND2_303(g14761,g12651,g10281);
  ND2 NAND2_304(I22844,g12113,g21228);
  ND4 NAND4_56(g21555,g17846,g14946,g17686,g17650);
  ND4 NAND4_57(g16854,g3965,g13824,g3976,g8595);
  ND2 NAND2_305(g11974,g2185,g8259);
  ND2 NAND2_306(g31671,I29262,I29263);
  ND4 NAND4_58(g27933,g21228,g25356,g26424,g26236);
  ND3 NAND3_49(g19549,g15969,g10841,g10899);
  ND4 NAND4_59(g8806,g358,g370,g376,g385);
  ND2 NAND2_307(g11639,g8933,g4722);
  ND2 NAND2_308(g9823,I13383,I13384);
  ND2 NAND2_309(g12933,g7150,g10515);
  ND2 NAND2_310(I25907,g26256,g24782);
  ND4 NAND4_60(g10207,g6315,g6358,g6329,g6351);
  ND2 NAND2_311(I20204,g16246,I20203);
  ND2 NAND2_312(g26752,g9397,g25189);
  ND2 NAND2_313(g14005,g11514,g11729);
  ND4 NAND4_61(g16660,g3953,g11225,g3969,g13933);
  ND2 NAND2_314(I26439,g26549,I26438);
  ND4 NAND4_62(g17605,g5559,g14425,g5630,g12563);
  ND2 NAND2_315(g11992,g7275,g1772);
  ND2 NAND2_316(I29314,g29501,I29313);
  ND2 NAND2_317(I26438,g26549,g14271);
  ND2 NAND2_318(I12096,g1339,g1322);
  ND2 NAND2_319(I23962,g23184,I23961);
  ND2 NAND2_320(I17446,g13336,g956);
  ND3 NAND3_50(g28206,g12546,g26105,g27985);
  ND2 NAND2_321(g25309,g22384,g12021);
  ND2 NAND2_322(I13564,g2648,g2652);
  ND2 NAND2_323(I12730,g4287,I12728);
  ND2 NAND2_324(g7857,I12241,I12242);
  ND3 NAND3_51(g28758,g27779,g7356,g7275);
  ND2 NAND2_325(I29269,g29486,g12050);
  ND4 NAND4_63(g14771,g5961,g12129,g5969,g12351);
  ND2 NAND2_326(g8913,I12877,I12878);
  ND3 NAND3_52(g11442,g8644,g3288,g3343);
  ND2 NAND2_327(I13183,g6500,I13182);
  ND2 NAND2_328(g14683,g12553,g12443);
  ND4 NAND4_64(g17514,g3917,g13772,g4019,g8595);
  ND2 NAND2_329(g25495,g12483,g22472);
  ND2 NAND2_330(g12592,I15364,I15365);
  ND2 NAND2_331(I13509,g2089,g2093);
  ND2 NAND2_332(I14247,g1322,g8091);
  ND2 NAND2_333(I15041,g9752,g1834);
  ND2 NAND2_334(g10515,g10337,g5022);
  ND2 NAND2_335(I13851,g862,I13850);
  ND2 NAND2_336(g25985,g24631,g23956);
  ND2 NAND2_337(g14882,g12558,g12453);
  ND2 NAND2_338(g34424,I32440,I32441);
  ND2 NAND2_339(g14407,g12008,g9807);
  ND3 NAND3_53(g19856,g13626,g16278,g8105);
  ND2 NAND2_340(I23951,g13603,I23949);
  ND2 NAND2_341(I15340,g10154,g2541);
  ND2 NAND2_342(g26255,g8075,g24779);
  ND2 NAND2_343(g12152,g2485,g8324);
  ND2 NAND2_344(g22325,g1252,g19140);
  ND2 NAND2_345(g13983,g11658,g8906);
  ND4 NAND4_65(g16694,g3905,g13772,g3976,g11631);
  ND4 NAND4_66(g17788,g5232,g14490,g5327,g12497);
  ND2 NAND2_346(g12413,g7521,g5654);
  ND2 NAND2_347(g10584,g7362,g7405);
  ND2 NAND2_348(g28406,g27064,g13675);
  ND2 NAND2_349(I13452,g1955,g1959);
  ND3 NAND3_54(g28962,g27886,g2040,g7369);
  ND2 NAND2_350(I29279,g12081,I29277);
  ND3 NAND3_55(g28500,g590,g27629,g12323);
  ND2 NAND2_351(g10759,g7537,g324);
  ND3 NAND3_56(g15721,g7564,g311,g13385);
  ND2 NAND2_352(I29278,g29488,I29277);
  ND2 NAND2_353(I14766,g5821,I14764);
  ND2 NAND2_354(I15130,g2527,I15128);
  ND2 NAND2_355(I15193,g9935,g6005);
  ND2 NAND2_356(I29286,g12085,I29284);
  ND2 NAND2_357(g14758,g7704,g12405);
  ND2 NAND2_358(g11130,g1221,g7918);
  ND2 NAND2_359(g14082,g11697,g11537);
  ND2 NAND2_360(g11193,I14258,I14259);
  ND3 NAND3_57(g13130,g1351,g11815,g11336);
  ND2 NAND2_361(g14107,g11571,g11527);
  ND3 NAND3_58(g16278,g8102,g8057,g13664);
  ND2 NAND2_362(g12020,g2028,g8365);
  ND3 NAND3_59(g19611,g1070,g1199,g15995);
  ND2 NAND2_363(g23139,g21163,g10756);
  ND3 NAND3_60(g16306,g4944,g13971,g12088);
  ND2 NAND2_364(I12261,g1454,g1448);
  ND2 NAND2_365(g14940,g12744,g12581);
  ND2 NAND2_366(I18627,g14712,I18625);
  ND3 NAND3_61(g13475,g1008,g11294,g11786);
  ND2 NAND2_367(g14848,g12651,g12453);
  ND4 NAND4_67(g27282,g11192,g26269,g26248,g479);
  ND4 NAND4_68(g21415,g17773,g14771,g17740,g14739);
  ND4 NAND4_69(g16815,g3909,g13824,g4005,g11631);
  ND4 NAND4_70(g13727,g174,g203,g168,g12812);
  ND4 NAND4_71(g15734,g5228,g12059,g5290,g14631);
  ND2 NAND2_368(g14804,g12651,g12798);
  ND2 NAND2_369(g25255,g20979,g23659);
  ND2 NAND2_370(I13731,g4537,I13729);
  ND2 NAND2_371(g12357,g7439,g6329);
  ND2 NAND2_372(g31978,g30580,g15591);
  ND2 NAND2_373(I22824,g21434,I22822);
  ND2 NAND2_374(I15253,g10078,g1848);
  ND2 NAND2_375(g24621,g22957,g2927);
  ND2 NAND2_376(I18681,g2638,I18680);
  ND2 NAND2_377(g14962,g12558,g10281);
  ND2 NAND2_378(g13600,g3021,g11039);
  ND2 NAND2_379(I22931,g21228,I22929);
  ND2 NAND2_380(g9645,g2060,g2028);
  ND2 NAND2_381(g23576,I22718,I22719);
  ND2 NAND2_382(g19764,I20166,I20167);
  ND2 NAND2_383(g11952,g1624,g8187);
  ND2 NAND2_384(I15175,g9977,I15174);
  ND2 NAND2_385(I32757,g34469,I32756);
  ND2 NAND2_386(I14370,g3303,I14368);
  ND2 NAND2_387(g26782,g9467,g25203);
  ND2 NAND2_388(g13821,g11251,g8340);
  ND2 NAND2_389(g14048,g11658,g11483);
  ND2 NAND2_390(I15264,g2273,I15262);
  ND2 NAND2_391(g22755,g20136,g18984);
  ND2 NAND2_392(g28421,g27074,g13715);
  ND3 NAND3_62(g26352,g744,g24875,g11679);
  ND2 NAND2_393(I12271,g956,I12269);
  ND3 NAND3_63(g13264,g11869,g11336,g11849);
  ND2 NAND2_394(g24933,g19466,g23154);
  ND4 NAND4_72(g13137,g10699,g7675,g1322,g1404);
  ND4 NAND4_73(g13516,g11533,g11490,g11444,g11412);
  ND2 NAND2_395(g15039,g12755,g7142);
  ND2 NAND2_396(g29060,g9649,g27800);
  ND4 NAND4_74(g17755,g5619,g14522,g5630,g9864);
  ND2 NAND2_397(g13873,g11566,g11729);
  ND2 NAND2_398(I31974,g33631,I31972);
  ND2 NAND2_399(g14947,g12785,g10491);
  ND2 NAND2_400(g10605,g2555,g7490);
  ND2 NAND2_401(g12482,I15307,I15308);
  ND3 NAND3_64(g25470,g22457,g2051,g8365);
  ND2 NAND2_402(g13834,g4754,g11773);
  ND3 NAND3_65(g16321,g4955,g13996,g12088);
  ND2 NAND2_403(g10951,g7845,g7868);
  ND3 NAND3_66(g28920,g27779,g1802,g7315);
  ND2 NAND2_404(g24574,g22709,g22687);
  ND2 NAND2_405(g14234,g9177,g11881);
  ND2 NAND2_406(g31706,I29270,I29271);
  ND2 NAND2_407(I18626,g2079,I18625);
  ND3 NAND3_67(g28946,g27907,g2495,g2421);
  ND2 NAND2_408(g25467,g12432,g22417);
  ND2 NAND2_409(g23761,I22893,I22894);
  ND2 NAND2_410(g23692,g9501,g20995);
  ND2 NAND2_411(g27380,I26071,I26072);
  ND2 NAND2_412(g12356,g7438,g6012);
  ND2 NAND2_413(g9591,g1926,g1894);
  ND3 NAND3_68(g12999,g4392,g10476,g4401);
  ND3 NAND3_69(g11320,g4633,g4621,g7202);
  ND2 NAND2_414(g25984,g24567,g22668);
  ND2 NAND2_415(g19886,g11403,g17794);
  ND2 NAND2_416(I15122,g9910,I15121);
  ND2 NAND2_417(g13346,g4854,g11012);
  ND2 NAND2_418(g19792,I20204,I20205);
  ND2 NAND2_419(I14957,g6181,I14955);
  ND3 NAND3_70(g26053,g22875,g24677,g22941);
  ND3 NAND3_71(g13464,g10831,g4793,g4776);
  ND2 NAND2_420(g13797,g8102,g11273);
  ND2 NAND2_421(g11292,I14331,I14332);
  ND2 NAND2_422(I32756,g34469,g25779);
  ND2 NAND2_423(g11153,I14205,I14206);
  ND2 NAND2_424(g29094,g27858,g9700);
  ND3 NAND3_72(g12449,g7004,g5297,g5352);
  ND2 NAND2_425(I14290,g8282,I14289);
  ND2 NAND2_426(g11409,g9842,g3298);
  ND2 NAND2_427(I22894,g21228,I22892);
  ND2 NAND2_428(I14427,g8595,g4005);
  ND4 NAND4_75(g14829,g6621,g12137,g6675,g12471);
  ND2 NAND2_429(I31983,g33653,g33648);
  ND2 NAND2_430(g14434,g6415,g11945);
  ND2 NAND2_431(g29018,g9586,g27742);
  ND2 NAND2_432(I12878,g4180,I12876);
  ND2 NAND2_433(g10946,g1489,g7876);
  ND3 NAND3_73(g28927,g27837,g1906,g7322);
  ND4 NAND4_76(g14946,g6247,g12173,g6346,g12672);
  ND2 NAND2_434(g9750,I13335,I13336);
  ND2 NAND2_435(I11826,g4601,I11824);
  ND2 NAND2_436(g14344,g5377,g11885);
  ND2 NAND2_437(g24583,g22753,g22711);
  ND2 NAND2_438(I13182,g6500,g6505);
  ND2 NAND2_439(I17496,g1448,I17494);
  ND3 NAND3_74(g28903,g27800,g2197,g7280);
  ND2 NAND2_440(g14682,g4933,g11780);
  ND2 NAND2_441(g12149,g8205,g2185);
  ND2 NAND2_442(I14481,g10074,I14480);
  ND3 NAND3_75(g28755,g27742,g7268,g1592);
  ND2 NAND2_443(g12148,g2060,g8310);
  ND4 NAND4_77(g13109,g6279,g12173,g6369,g10003);
  ND4 NAND4_78(g16772,g3558,g13799,g3654,g11576);
  ND2 NAND2_444(g24787,g3391,g23079);
  ND3 NAND3_76(g29001,g27937,g2599,g7431);
  ND4 NAND4_79(g13108,g5551,g12029,g5685,g9864);
  ND2 NAND2_445(g12343,g7470,g5630);
  ND3 NAND3_77(g13283,g12440,g12399,g9843);
  ND2 NAND2_446(I22801,g21434,I22799);
  ND3 NAND3_78(g11492,g6928,g6941,g8756);
  ND3 NAND3_79(g12971,g9024,g8977,g10664);
  ND2 NAND2_447(I12545,g191,I12544);
  ND2 NAND2_448(g9528,I13183,I13184);
  ND2 NAND2_449(g12369,g9049,g637);
  ND2 NAND2_450(g28395,g27074,g13655);
  ND2 NAND2_451(I14956,g9620,I14955);
  ND2 NAND2_452(g11381,g9660,g3274);
  ND2 NAND2_453(g28899,g27833,g14612);
  ND2 NAND2_454(I18529,g1811,g14640);
  ND2 NAND2_455(g28990,g27882,g8310);
  ND3 NAND3_80(g17220,g9369,g9298,g14376);
  ND2 NAND2_456(I15174,g9977,g2661);
  ND2 NAND2_457(g29157,g9835,g27937);
  ND3 NAND3_81(g17246,g9439,g9379,g14405);
  ND3 NAND3_82(g12412,g10044,g5297,g5348);
  ND2 NAND2_458(I26049,g25997,g13500);
  ND3 NAND3_83(g26382,g577,g24953,g12323);
  ND3 NAND3_84(g33930,g33394,g12767,g9848);
  ND2 NAND2_459(g22754,g20114,g19376);
  ND2 NAND2_460(g33838,g33083,g4369);
  ND2 NAND2_461(g14927,g12695,g10281);
  ND2 NAND2_462(g16586,g13851,g13823);
  ND2 NAND2_463(I22866,g21228,I22864);
  ND2 NAND2_464(g21345,g11429,g17157);
  ND3 NAND3_85(g27582,g10857,g26131,g26105);
  ND2 NAND2_465(g9372,g5080,g5084);
  ND3 NAND3_86(g28861,g27837,g7405,g1906);
  ND2 NAND2_466(I20461,g17515,I20460);
  ND3 NAND3_87(g25476,g22472,g2476,g8373);
  ND2 NAND2_467(g8359,I12545,I12546);
  ND2 NAND2_468(g24662,g22957,g2955);
  ND2 NAND2_469(I24461,g23796,g14437);
  ND2 NAND2_470(g10604,g7424,g7456);
  ND4 NAND4_80(g15751,g5591,g14522,g5666,g14669);
  ND4 NAND4_81(g10755,g7352,g7675,g1322,g1404);
  ND2 NAND2_471(g24890,g13852,g22929);
  ND2 NAND2_472(g14755,g12593,g12772);
  ND3 NAND3_88(g19495,g15969,g10841,g7781);
  ND2 NAND2_473(g27925,I26439,I26440);
  ND2 NAND2_474(I22923,g21284,I22921);
  ND2 NAND2_475(g29660,g28448,g9582);
  ND3 NAND3_89(g20248,g17056,g14146,g14123);
  ND2 NAND2_476(g16275,g9291,g13480);
  ND2 NAND2_477(g14981,g12785,g12632);
  ND2 NAND2_478(I14211,g9252,g9295);
  ND2 NAND2_479(g9334,g827,g832);
  ND2 NAND2_480(g12112,g8139,g1624);
  ND2 NAND2_481(I17923,g13378,g1478);
  ND3 NAND3_90(g33306,g776,g32212,g11679);
  ND4 NAND4_82(g11326,g8993,g376,g365,g370);
  ND2 NAND2_482(g20081,g11325,g17794);
  ND2 NAND2_483(g14794,g12492,g12772);
  ND2 NAND2_484(g14845,g12558,g12798);
  ND2 NAND2_485(I14497,g9020,g8737);
  ND2 NAND2_486(I24365,g14320,I24363);
  ND2 NAND2_487(I13850,g862,g7397);
  ND4 NAND4_83(g13040,g5196,g12002,g5308,g9780);
  ND2 NAND2_488(g13948,g11610,g8864);
  ND2 NAND2_489(g14899,g12744,g10421);
  ND2 NAND2_490(g29085,g9694,g27837);
  ND2 NAND2_491(g28997,g27903,g8324);
  ND2 NAND2_492(g25382,g12333,g22342);
  ND2 NAND2_493(I12289,g1300,I12287);
  ND4 NAND4_84(g14898,g5901,g12129,g6000,g12614);
  ND2 NAND2_494(I32204,g33670,I32202);
  ND2 NAND2_495(I23950,g23162,I23949);
  ND2 NAND2_496(g15014,g12785,g12680);
  ND2 NAND2_497(I12288,g1484,I12287);
  ND2 NAND2_498(g24380,I23601,I23602);
  ND2 NAND2_499(g12429,g7473,g6675);
  ND2 NAND2_500(g14521,g12170,g5428);
  ND2 NAND2_501(I25221,g24718,I25219);
  ND2 NAND2_502(g12428,g7472,g6358);
  ND3 NAND3_91(g28871,g27858,g7418,g2331);
  ND2 NAND2_503(I17885,g1135,I17883);
  ND2 NAND2_504(g9908,I13453,I13454);
  ND2 NAND2_505(g22902,g18957,g2848);
  ND2 NAND2_506(I16780,g12332,I16778);
  ND2 NAND2_507(g10573,g7992,g8179);
  ND2 NAND2_508(g9567,g6116,g6120);
  ND2 NAND2_509(g14861,g12744,g10341);
  ND2 NAND2_510(g14573,g9506,g12249);
  ND2 NAND2_511(g24932,g19886,g23172);
  ND4 NAND4_85(g15720,g5917,g14497,g6019,g9935);
  ND3 NAND3_92(g11933,g837,g9334,g7197);
  ND2 NAND2_512(I14855,g5142,I14853);
  ND2 NAND2_513(g14045,g11571,g11747);
  ND2 NAND2_514(g29335,g25540,g28131);
  ND2 NAND2_515(g13634,g11797,g11261);
  ND2 NAND2_516(g13851,g8224,g11360);
  ND2 NAND2_517(g27317,g24793,g26255);
  ND2 NAND2_518(I12374,g3462,I12372);
  ND2 NAND2_519(g25215,I24384,I24385);
  ND2 NAND2_520(g7850,g554,g807);
  ND2 NAND2_521(g12317,g10026,g6486);
  ND2 NAND2_522(g29694,g28391,g13709);
  ND2 NAND2_523(g14098,g11566,g8864);
  ND2 NAND2_524(g17699,I18681,I18682);
  ND2 NAND2_525(g25439,g22498,g12122);
  ND3 NAND3_93(g28911,g27907,g7456,g2465);
  ND2 NAND2_526(g23972,g7097,g20751);
  ND3 NAND3_94(g17290,g9506,g9449,g14431);
  ND2 NAND2_527(I29253,g29482,g12017);
  ND2 NAND2_528(g29131,g27907,g9762);
  ND2 NAND2_529(I15213,g10035,I15212);
  ND2 NAND2_530(I12842,g4235,I12840);
  ND2 NAND2_531(g25349,g22432,g12051);
  ND2 NAND2_532(g12245,g7344,g5637);
  ND2 NAND2_533(g12323,g9480,g640);
  ND2 NAND2_534(I14714,g5128,I14712);
  ND2 NAND2_535(g22661,g20136,g94);
  ND2 NAND2_536(I13730,g4534,I13729);
  ND4 NAND4_86(g27775,g21228,g25262,g26424,g26166);
  ND3 NAND3_95(g16236,g13573,g13554,g13058);
  ND2 NAND2_537(I14257,g8154,g3133);
  ND3 NAND3_96(g28950,g27937,g7490,g2599);
  ND2 NAND2_538(I15051,g9759,g2259);
  ND2 NAND2_539(I14818,g6513,I14816);
  ND2 NAND2_540(g9724,g5092,g5084);
  ND2 NAND2_541(g22715,g20114,g2999);
  ND2 NAND2_542(I23120,g417,I23118);
  ND2 NAND2_543(g24620,g22902,g22874);
  ND4 NAND4_87(g14871,g6653,g12211,g6661,g12471);
  ND2 NAND2_544(I12544,g191,g194);
  ND2 NAND2_545(g13756,g203,g12812);
  ND2 NAND2_546(I18680,g2638,g14752);
  ND2 NAND2_547(g12232,g8804,g4878);
  ND3 NAND3_97(g16264,g518,g9158,g13223);
  ND2 NAND2_548(g19875,g13667,g16316);
  ND2 NAND2_549(I22930,g12223,I22929);
  ND3 NAND3_98(g26052,g22714,g24662,g22921);
  ND2 NAND2_550(g26745,g6856,g25317);
  ND4 NAND4_88(g17572,g3598,g13799,g3676,g8542);
  ND2 NAND2_551(g11350,I14369,I14370);
  ND2 NAND2_552(I22965,g12288,g21228);
  ND2 NAND2_553(I32433,g34051,I32431);
  ND2 NAND2_554(g24369,I23586,I23587);
  ND2 NAND2_555(g12512,g7766,g10312);
  ND2 NAND2_556(g21359,g11509,g17157);
  ND2 NAND2_557(g13846,g1116,g10649);
  ND2 NAND2_558(g10472,I13851,I13852);
  ND2 NAND2_559(g11396,g8713,g4688);
  ND2 NAND2_560(I12270,g1141,I12269);
  ND2 NAND2_561(I14735,g5475,I14733);
  ND3 NAND3_99(g19455,g15969,g10841,g7781);
  ND4 NAND4_89(g20133,g17668,g17634,g17597,g14569);
  ND2 NAND2_562(g17297,g2729,g14291);
  ND2 NAND2_563(g21344,g11428,g17157);
  ND4 NAND4_90(g11405,g2741,g2735,g6856,g2748);
  ND4 NAND4_91(g15781,g6267,g12173,g6329,g14745);
  ND2 NAND2_564(g20011,g3731,g16476);
  ND2 NAND2_565(g14776,g12780,g12622);
  ND3 NAND3_100(g28203,g12546,g27985,g27977);
  ND3 NAND3_101(g10754,g7936,g7913,g8411);
  ND2 NAND2_566(g29015,g27742,g9586);
  ND2 NAND2_567(g13929,g11669,g11763);
  ND2 NAND2_568(I12219,g1478,I12217);
  ND2 NAND2_569(g25200,g5742,g23642);
  ND2 NAND2_570(g14825,g12806,g12680);
  ND2 NAND2_571(g14950,g7812,g12632);
  ND2 NAND2_572(g11020,g9187,g9040);
  ND2 NAND2_573(g12080,g1917,g8201);
  ND4 NAND4_92(g13928,g3562,g11238,g3680,g11576);
  ND2 NAND2_574(I12218,g1437,I12217);
  ND2 NAND2_575(g14858,g7766,g12515);
  ND2 NAND2_576(g19782,I20188,I20189);
  ND2 NAND2_577(g29556,g28349,g13486);
  ND2 NAND2_578(g31747,I29296,I29297);
  ND2 NAND2_579(g14151,g11692,g11483);
  ND2 NAND2_580(g14996,g12662,g10312);
  ND2 NAND2_581(g24925,g20092,g23154);
  ND2 NAND2_582(g24958,g21330,g23462);
  ND4 NAND4_93(g17520,g5260,g12002,g5276,g14631);
  ND2 NAND2_583(g12461,g7536,g6000);
  ND2 NAND2_584(I24364,g23687,I24363);
  ND3 NAND3_102(g12342,g7004,g7018,g10129);
  ND2 NAND2_585(I22937,g12226,I22936);
  ND2 NAND2_586(I26395,g14227,I26393);
  ND2 NAND2_587(I14923,g9558,g5835);
  ND2 NAND2_588(g12145,g8195,g1760);
  ND2 NAND2_589(g11302,g9496,g3281);
  ND2 NAND2_590(I15105,g9780,g5313);
  ND2 NAND2_591(I23980,g13670,I23978);
  ND2 NAND2_592(g24944,g21354,g23363);
  ND4 NAND4_94(g13105,g10671,g7675,g1322,g1404);
  ND2 NAND2_593(I16779,g11292,I16778);
  ND2 NAND2_594(I12470,g392,I12468);
  ND2 NAND2_595(g9092,g3004,g3050);
  ND2 NAND2_596(I16778,g11292,g12332);
  ND3 NAND3_103(g19589,g15969,g10841,g10884);
  ND2 NAND2_597(I12277,g1467,g1472);
  ND2 NAND2_598(I13499,g232,I13497);
  ND2 NAND2_599(I17884,g13336,I17883);
  ND2 NAND2_600(g15021,g12711,g10341);
  ND2 NAND2_601(I12075,g996,I12074);
  ND2 NAND2_602(g27365,I26050,I26051);
  ND2 NAND2_603(g24802,I23970,I23971);
  ND2 NAND2_604(g29186,g27051,g4507);
  ND2 NAND2_605(g29676,g28381,g13676);
  ND3 NAND3_104(g7690,g4669,g4659,g4653);
  ND4 NAND4_95(g15726,g6263,g14529,g6365,g10003);
  ND2 NAND2_606(I13498,g255,I13497);
  ND2 NAND2_607(g24793,g3742,g23124);
  ND2 NAND2_608(g26235,g8016,g24766);
  ND2 NAND2_609(g14058,g7121,g11537);
  ND2 NAND2_610(I26440,g14271,I26438);
  ND2 NAND2_611(g28895,g27775,g8146);
  ND2 NAND2_612(I14885,g5489,I14883);
  ND2 NAND2_613(g11881,g9060,g3361);
  ND2 NAND2_614(I14854,g9433,I14853);
  ND2 NAND2_615(g25400,g22472,g12086);
  ND2 NAND2_616(g12225,g8324,g2453);
  ND2 NAND2_617(g14902,g7791,g12581);
  ND2 NAND2_618(g12471,I15288,I15289);
  ND2 NAND2_619(I29303,g29496,I29302);
  ND2 NAND2_620(g12087,g7431,g2599);
  ND2 NAND2_621(g14120,g11780,g4907);
  ND4 NAND4_96(g14739,g5929,g12067,g5983,g12351);
  ND2 NAND2_622(g10738,g6961,g10308);
  ND2 NAND2_623(I22922,g14677,I22921);
  ND2 NAND2_624(I25845,g26212,g24799);
  ND2 NAND2_625(g14146,g11020,g691);
  ND2 NAND2_626(g32072,g31009,g13301);
  ND2 NAND2_627(g19466,g11562,g17794);
  ND2 NAND2_628(I15003,g9691,I15002);
  ND2 NAND2_629(g12244,g7343,g5320);
  ND3 NAND3_105(g13248,g9985,g12399,g9843);
  ND2 NAND2_630(I14480,g10074,g655);
  ND2 NAND2_631(g28376,g27064,g13620);
  ND2 NAND2_632(g13779,g11804,g11283);
  ND2 NAND2_633(I22685,g21434,I22683);
  ND2 NAND2_634(g27955,I26460,I26461);
  ND2 NAND2_635(g28980,g27933,g14680);
  ND2 NAND2_636(I23987,g482,I23985);
  ND2 NAND2_637(g23719,I22845,I22846);
  ND2 NAND2_638(I12401,g3808,g3813);
  ND2 NAND2_639(g28888,g27738,g8139);
  ND3 NAND3_106(g28824,g27779,g7356,g1772);
  ND2 NAND2_640(I20488,g16757,I20486);
  ND2 NAND2_641(I22800,g11960,I22799);
  ND2 NAND2_642(I22936,g12226,g21228);
  ND2 NAND2_643(g11356,g9552,g3632);
  ND4 NAND4_97(g8691,g3267,g3310,g3281,g3303);
  ND2 NAND2_644(g13945,g691,g11740);
  ND3 NAND3_107(g19874,g13665,g16299,g8163);
  ND4 NAND4_98(g17581,g5607,g12029,g5623,g14669);
  ND3 NAND3_108(g17315,g9564,g9516,g14503);
  ND3 NAND3_109(g28931,g27886,g2070,g1996);
  ND2 NAND2_645(I23969,g22202,g490);
  ND2 NAND2_646(g14547,g9439,g12201);
  ND2 NAND2_647(g14895,g7766,g12571);
  ND2 NAND2_648(g11998,g8324,g8373);
  ND2 NAND2_649(I22762,g21434,I22760);
  ND2 NAND2_650(g13672,g8933,g11261);
  ND2 NAND2_651(g12459,g7437,g5623);
  ND4 NAND4_99(g16663,g13854,g13834,g14655,g12292);
  ND2 NAND2_652(g10551,g1728,g7356);
  ND2 NAND2_653(g21388,g11608,g17157);
  ND3 NAND3_110(g24880,g23281,g23266,g22839);
  ND2 NAND2_654(g23324,g703,g20181);
  ND2 NAND2_655(g14572,g12169,g9678);
  ND2 NAND2_656(I14734,g9732,I14733);
  ND2 NAND2_657(I20189,g1333,I20187);
  ND2 NAND2_658(g21272,g11268,g17157);
  ND2 NAND2_659(I13043,g5115,g5120);
  ND2 NAND2_660(I14993,g6527,I14991);
  ND2 NAND2_661(I20188,g16272,I20187);
  ND3 NAND3_111(g13513,g1351,g11815,g8002);
  ND2 NAND2_662(g14127,g11653,g11435);
  ND4 NAND4_100(g21462,g17816,g14871,g17779,g14829);
  ND2 NAND2_663(g11961,g9777,g5105);
  ND2 NAND2_664(g12079,g1792,g8195);
  ND2 NAND2_665(g28860,g27775,g14586);
  ND4 NAND4_101(g13897,g3211,g11217,g3329,g11519);
  ND2 NAND2_666(I20460,g17515,g14187);
  ND2 NAND2_667(I24383,g23721,g14347);
  ND2 NAND2_668(g12078,g8187,g8093);
  ND2 NAND2_669(I26071,g26026,I26070);
  ND2 NAND2_670(I15212,g10035,g1714);
  ND2 NAND2_671(g14956,g12604,g10281);
  ND2 NAND2_672(I11879,g4430,I11877);
  ND2 NAND2_673(g14889,g12609,g12824);
  ND4 NAND4_102(g16757,g13911,g13886,g14120,g11675);
  ND2 NAND2_674(I11878,g4388,I11877);
  ND3 NAND3_112(g28987,g27886,g2070,g7411);
  ND3 NAND3_113(g25435,g22432,g2342,g8316);
  ND2 NAND2_675(I23979,g23198,I23978);
  ND2 NAND2_676(g24989,g21345,g23363);
  ND2 NAND2_677(g12159,g8765,g4864);
  ND2 NAND2_678(g12125,g9728,g5101);
  ND2 NAND2_679(I21978,g19620,I21976);
  ND2 NAND2_680(I22974,g19638,I22972);
  ND2 NAND2_681(I23978,g23198,g13670);
  ND2 NAND2_682(g24988,g546,g23088);
  ND2 NAND2_683(g24924,g20007,g23172);
  ND2 NAND2_684(I15149,g5659,I15147);
  ND2 NAND2_685(g21360,g11510,g17157);
  ND2 NAND2_686(I23986,g22182,I23985);
  ND2 NAND2_687(g27295,g24776,g26208);
  ND4 NAND4_103(g20271,g16925,g14054,g16657,g16628);
  ND2 NAND2_688(g11149,g1564,g7948);
  ND2 NAND2_689(I15148,g9864,I15147);
  ND2 NAND2_690(g28969,g27854,g8267);
  ND2 NAND2_691(I26367,g26400,I26366);
  ND2 NAND2_692(I26394,g26488,I26393);
  ND2 NAND2_693(g12144,I15003,I15004);
  ND2 NAND2_694(g9543,g2217,g2185);
  ND4 NAND4_104(g13097,g5204,g12002,g5339,g9780);
  ND2 NAND2_695(g10520,g7195,g7115);
  ND2 NAND2_696(g13104,g1404,g10794);
  ND2 NAND2_697(g12336,I15175,I15176);
  ND2 NAND2_698(g14520,g9369,g12163);
  ND2 NAND2_699(I14187,g3470,I14185);
  ND2 NAND2_700(g7150,g5016,g5062);
  ND2 NAND2_701(I25220,g482,I25219);
  ND4 NAND4_105(g20199,g16815,g13968,g16749,g13907);
  ND2 NAND2_702(g11971,g8249,g8302);
  ND2 NAND2_703(g28870,g27796,g14588);
  ND3 NAND3_114(g34048,g33669,g10583,g7442);
  ND2 NAND2_704(I13079,g5467,I13077);
  ND2 NAND2_705(I13444,g239,I13442);
  ND2 NAND2_706(I32432,g34056,I32431);
  ND2 NAND2_707(g14546,g12125,g9613);
  ND2 NAND2_708(g14089,g11755,g4717);
  ND2 NAND2_709(g22688,g20219,g2936);
  ND4 NAND4_106(g20198,g16813,g13958,g16745,g13927);
  ND4 NAND4_107(g17706,g3921,g11255,g3983,g13933);
  ND4 NAND4_108(g17597,g3191,g13700,g3303,g8481);
  ND2 NAND2_710(I12074,g996,g979);
  ND2 NAND2_711(I13078,g5462,I13077);
  ND4 NAND4_109(g14088,g3901,g11255,g4000,g11631);
  ND2 NAND2_712(g14024,g7121,g11763);
  ND4 NAND4_110(g17689,g6645,g12137,g6661,g14786);
  ND2 NAND2_713(I18589,g14679,I18587);
  ND2 NAND2_714(g24528,g4098,g22654);
  ND2 NAND2_715(g17624,I18588,I18589);
  ND3 NAND3_115(g28867,g27800,g2227,g2153);
  ND2 NAND2_716(I18588,g2370,I18587);
  ND2 NAND2_717(g7836,g4653,g4688);
  ND2 NAND2_718(I20467,g16663,g16728);
  ND2 NAND2_719(I14169,g8389,g3119);
  ND2 NAND2_720(I14884,g9500,I14883);
  ND3 NAND3_116(g11412,g8666,g6918,g8697);
  ND2 NAND2_721(g15702,g13066,g7293);
  ND2 NAND2_722(g13850,g11279,g8396);
  ND2 NAND2_723(g15904,I17380,I17381);
  ND2 NAND2_724(g25049,g21344,g23462);
  ND3 NAND3_117(g12289,g9978,g9766,g9708);
  ND2 NAND2_725(g14659,g12646,g12443);
  ND4 NAND4_111(g14625,g3897,g11225,g4031,g8595);
  ND4 NAND4_112(g14987,g6593,g12211,g6692,g12721);
  ND4 NAND4_113(g20161,g17732,g17706,g17670,g14625);
  ND2 NAND2_726(g22885,g9104,g20154);
  ND2 NAND2_727(g12023,g2453,g8373);
  ND2 NAND2_728(g28910,g27854,g14614);
  ND4 NAND4_114(g13896,g3227,g11194,g3281,g11350);
  ND2 NAND2_729(I23917,g23975,g9333);
  ND2 NAND2_730(g25048,g542,g23088);
  ND2 NAND2_731(g12224,I15088,I15089);
  ND2 NAND2_732(g14943,g7791,g12622);
  ND2 NAND2_733(I13336,g1691,I13334);
  ND2 NAND2_734(g27687,g25200,g26714);
  ND2 NAND2_735(g14968,g12739,g10312);
  ND2 NAND2_736(g11959,g8316,g2342);
  ND2 NAND2_737(g13627,g11172,g8388);
  ND2 NAND2_738(I22684,g11893,I22683);
  ND2 NAND2_739(I20167,g990,I20165);
  ND2 NAND2_740(g14855,g12700,g12824);
  ND2 NAND2_741(I12729,g4291,I12728);
  ND4 NAND4_115(g13050,g5543,g12029,g5654,g9864);
  ND4 NAND4_116(g13958,g3610,g11238,g3618,g11389);
  ND2 NAND2_742(I12728,g4291,g4287);
  ND3 NAND3_118(g28877,g27937,g7490,g7431);
  ND2 NAND2_743(g20068,g11293,g17794);
  ND2 NAND2_744(I26366,g26400,g14211);
  ND2 NAND2_745(I14531,g8840,I14530);
  ND2 NAND2_746(g13742,g11780,g11283);
  ND2 NAND2_747(g11944,I14765,I14766);
  ND2 NAND2_748(g7620,I12097,I12098);
  ND2 NAND2_749(g8010,I12345,I12346);
  ND2 NAND2_750(I14186,g8442,I14185);
  ND2 NAND2_751(g17287,g7262,g14228);
  ND2 NAND2_752(g12195,g2619,g8381);
  ND2 NAND2_753(g17596,g8686,g14367);
  ND2 NAND2_754(g25514,g12540,g22498);
  ND2 NAND2_755(g24792,I23950,I23951);
  ND2 NAND2_756(g17243,g7247,g14212);
  ND2 NAND2_757(g12525,g7522,g6668);
  ND2 NAND2_758(g12016,g1648,g8093);
  ND2 NAND2_759(g23281,g18957,g2898);
  ND2 NAND2_760(g21301,g11371,g17157);
  ND2 NAND2_761(g21377,g11560,g17157);
  ND2 NAND2_762(g14055,g11697,g11763);
  ND4 NAND4_117(g17773,g5965,g14549,g5976,g9935);
  ND2 NAND2_763(I18485,g1677,g14611);
  ND2 NAND2_764(g14978,g12716,g10491);
  ND4 NAND4_118(g15780,g5937,g14549,g6012,g14701);
  ND2 NAND2_765(I17475,g13336,I17474);
  ND4 NAND4_119(g14590,g3546,g11207,g3680,g8542);
  ND2 NAND2_766(g24918,g136,g23088);
  ND4 NAND4_120(g17670,g3893,g13772,g4005,g8595);
  ND2 NAND2_767(g22839,g20114,g2988);
  ND2 NAND2_768(g23699,g21012,g11160);
  ND2 NAND2_769(I29302,g29496,g12121);
  ND2 NAND2_770(g25473,g12437,g22432);
  ND2 NAND2_771(g14741,g12711,g10421);
  ND2 NAND2_772(g27705,g25237,g26782);
  ND2 NAND2_773(g22838,g20219,g2960);
  ND4 NAND4_121(g17734,g5272,g14490,g5283,g9780);
  ND2 NAND2_774(g28923,g27775,g8195);
  ND3 NAND3_119(g16282,g4933,g13939,g12088);
  ND2 NAND2_775(g9442,g5424,g5428);
  ND2 NAND2_776(g27679,g25186,g26685);
  ND2 NAND2_777(I15129,g9914,I15128);
  ND2 NAND2_778(g12042,g9086,g703);
  ND2 NAND2_779(I15002,g9691,g1700);
  ND2 NAND2_780(I26095,g13539,I26093);
  ND2 NAND2_781(g12255,g9958,g6140);
  ND2 NAND2_782(g11002,g7475,g862);
  ND2 NAND2_783(I15128,g9914,g2527);
  ND2 NAND2_784(g13057,g969,g11294);
  ND2 NAND2_785(g14735,g12739,g12571);
  ND2 NAND2_786(g12188,g8249,g1894);
  ND2 NAND2_787(g12124,g8741,g4674);
  ND2 NAND2_788(I13392,g1825,I13390);
  ND3 NAND3_120(g11245,g7636,g7733,g7697);
  ND2 NAND2_789(I15299,g10112,I15298);
  ND3 NAND3_121(g12460,g10093,g5644,g5694);
  ND3 NAND3_122(g12686,g7097,g6682,g6736);
  ND2 NAND2_790(I20166,g16246,I20165);
  ND2 NAND2_791(g11323,I14351,I14352);
  ND4 NAND4_122(g14695,g5583,g12029,g5637,g12301);
  ND2 NAND2_792(g14018,g10323,g11483);
  ND2 NAND2_793(I15298,g10112,g1982);
  ND3 NAND3_123(g11533,g6905,g3639,g3698);
  ND2 NAND2_794(g21403,g11652,g17157);
  ND2 NAND2_795(g20783,g14616,g17225);
  ND3 NAND3_124(g12294,g10044,g7018,g10090);
  ND2 NAND2_796(g17618,I18580,I18581);
  ND3 NAND3_125(g28885,g27742,g1668,g7268);
  ND4 NAND4_123(g22306,g4584,g4616,g13202,g19071);
  ND2 NAND2_797(I22873,g21228,I22871);
  ND2 NAND2_798(I11865,g4434,I11864);
  ND2 NAND2_799(I14230,g8055,I14228);
  ND4 NAND4_124(g17468,g3215,g13700,g3317,g8481);
  ND2 NAND2_800(I21993,g7670,I21992);
  ND4 NAND4_125(g15787,g6283,g14575,g6358,g14745);
  ND4 NAND4_126(g14706,g6287,g12101,g6369,g12672);
  ND2 NAND2_801(I14992,g9685,I14991);
  ND4 NAND4_127(g21385,g17736,g14696,g17679,g14636);
  ND2 NAND2_802(I14510,g8721,I14508);
  ND4 NAND4_128(g15743,g5893,g14497,g6005,g9935);
  ND2 NAND2_803(g21354,g11468,g17157);
  ND2 NAND2_804(g14688,g12604,g12453);
  ND3 NAND3_126(g28287,g10504,g26131,g26973);
  ND2 NAND2_805(g12915,g12806,g12632);
  ND2 NAND2_806(I13383,g269,I13382);
  ND2 NAND2_807(g11445,g9771,g3976);
  ND2 NAND2_808(g14157,g11715,g11763);
  ND2 NAND2_809(g22666,g18957,g2878);
  ND4 NAND4_129(g13499,g11479,g11442,g11410,g11382);
  ND2 NAND2_810(I13065,g4308,g4304);
  ND2 NAND2_811(g14066,g11514,g11473);
  ND4 NAND4_130(g13498,g12577,g12522,g12462,g12416);
  ND2 NAND2_812(I15080,g1968,I15078);
  ND2 NAND2_813(g17363,g8635,g14367);
  ND3 NAND3_127(g28942,g27858,g2331,g7335);
  ND2 NAND2_814(g17217,g7239,g14194);
  ND2 NAND2_815(g21190,g6077,g17420);
  ND2 NAND2_816(g14876,g12492,g12443);
  ND2 NAND2_817(g14885,g12651,g12505);
  ND4 NAND4_131(g14854,g5555,g12093,g5654,g12563);
  ND3 NAND3_128(g10511,g4628,g7202,g4621);
  ND2 NAND2_818(g11432,g10295,g8864);
  ND2 NAND2_819(I23601,g22360,I23600);
  ND2 NAND2_820(g13432,g4793,g10831);
  ND2 NAND2_821(I14275,g8218,g3484);
  ND2 NAND2_822(g12155,g7753,g7717);
  ND4 NAND4_132(g12822,g6978,g7236,g7224,g7163);
  ND2 NAND2_823(g15027,g12667,g10341);
  ND2 NAND2_824(I15342,g2541,I15340);
  ND2 NAND2_825(g28930,g27833,g8201);
  ND2 NAND2_826(I24439,g23771,I24438);
  ND2 NAND2_827(g28965,g27882,g8255);
  ND2 NAND2_828(g30573,g29355,g19666);
  ND2 NAND2_829(I24438,g23771,g14411);
  ND2 NAND2_830(g15710,g319,g13385);
  ND2 NAND2_831(g9715,g5011,g4836);
  ND2 NAND2_832(g28131,g27051,g25838);
  ND3 NAND3_129(g31509,g599,g29933,g12323);
  ND2 NAND2_833(g10916,g1146,g7854);
  ND2 NAND2_834(I12241,g1111,I12240);
  ND4 NAND4_133(g33933,g33394,g12491,g12819,g12796);
  ND2 NAND2_835(g12589,g7591,g6692);
  ND2 NAND2_836(g12194,g8373,g8273);
  ND2 NAND2_837(g10550,g7268,g7308);
  ND4 NAND4_134(g13529,g11590,g11544,g11492,g11446);
  ND2 NAND2_838(I14517,g10147,I14516);
  ND3 NAND3_130(g12588,g10169,g6336,g6386);
  ND2 NAND2_839(g27401,I26094,I26095);
  ND3 NAND3_131(g12524,g7074,g7087,g10212);
  ND2 NAND2_840(g23659,g9434,g20854);
  ND2 NAND2_841(g11330,g9483,g1193);
  ND3 NAND3_132(g13528,g11294,g7549,g1008);
  ND2 NAND2_842(g13330,g4664,g11006);
  ND2 NAND2_843(g10307,I13730,I13731);
  ND2 NAND2_844(I15365,g2675,I15363);
  ND2 NAND2_845(g14085,g7121,g11584);
  ND4 NAND4_135(g17740,g5945,g14497,g6012,g12351);
  ND2 NAND2_846(g13764,g11252,g3072);
  ND2 NAND2_847(g8238,I12469,I12470);
  ND4 NAND4_136(g14596,g12196,g9775,g12124,g9663);
  ND2 NAND2_848(g12119,g2351,g8267);
  ND4 NAND4_137(g14054,g3550,g11238,g3649,g11576);
  ND2 NAND2_849(I22711,g11915,I22710);
  ND3 NAND3_133(g7701,g4859,g4849,g4843);
  ND4 NAND4_138(g21339,g15725,g13084,g15713,g13050);
  ND2 NAND2_850(g13960,g11669,g11537);
  ND2 NAND2_851(g32057,g31003,g13297);
  ND2 NAND2_852(g12118,g8259,g8150);
  ND2 NAND2_853(g12022,g7335,g2331);
  ND4 NAND4_139(g21338,g15741,g15734,g15728,g13097);
  ND2 NAND2_854(I26070,g26026,g13517);
  ND2 NAND2_855(I17474,g13336,g1105);
  ND4 NAND4_140(g16723,g3606,g13730,g3676,g11576);
  ND2 NAND2_856(g14773,g12711,g12581);
  ND3 NAND3_134(g24544,g22666,g22661,g22651);
  ND2 NAND2_857(g13709,g11755,g11261);
  ND2 NAND2_858(g25389,g22457,g12082);
  ND2 NAND2_859(g12285,I15122,I15123);
  ND2 NAND2_860(I15087,g9832,g2393);
  ND2 NAND2_861(g14655,g4743,g11755);
  ND2 NAND2_862(g11708,g10147,g10110);
  ND2 NAND2_863(g13708,g11200,g8507);
  ND2 NAND2_864(g12053,g2587,g8418);
  ND2 NAND2_865(g16097,g13319,g10998);
  ND2 NAND2_866(I26094,g26055,I26093);
  ND2 NAND2_867(I24415,g23751,I24414);
  ND2 NAND2_868(I15043,g1834,I15041);
  ND2 NAND2_869(g13043,g10521,g969);
  ND2 NAND2_870(g14930,g12609,g12515);
  ND2 NAND2_871(g14993,g12695,g12453);
  ND2 NAND2_872(I17381,g1129,I17379);
  ND2 NAND2_873(g24678,g22994,g23010);
  ND2 NAND2_874(g14838,g12492,g12405);
  ND2 NAND2_875(g14965,g12609,g12571);
  ND2 NAND2_876(g22908,g9104,g20175);
  ND4 NAND4_141(g13069,g5889,g12067,g6000,g9935);
  ND2 NAND2_877(g29702,g28395,g13712);
  ND3 NAND3_135(g34162,g785,g33823,g11679);
  ND2 NAND2_878(g15717,g10754,g13092);
  ND2 NAND2_879(I13401,g2246,g2250);
  ND2 NAND2_880(g11955,g8302,g1917);
  ND2 NAND2_881(g13955,g11621,g11527);
  ND2 NAND2_882(g11970,g1760,g8241);
  ND2 NAND2_883(g28410,g27074,g13679);
  ND2 NAND2_884(g19962,g11470,g17794);
  ND2 NAND2_885(g10618,g10153,g9913);
  ND2 NAND2_886(I14351,g8890,I14350);
  ND2 NAND2_887(g27693,g25216,g26752);
  ND2 NAND2_888(I11864,g4434,g4401);
  ND2 NAND2_889(g34220,I32186,I32187);
  ND2 NAND2_890(g28363,g27064,g13593);
  ND2 NAND2_891(g17568,I18486,I18487);
  ND2 NAND2_892(g14279,g12111,g9246);
  ND2 NAND2_893(g7887,I12278,I12279);
  ND2 NAND2_894(I13749,g4608,g4584);
  ND2 NAND2_895(g13886,g11804,g4922);
  ND2 NAND2_896(g7228,g6398,g6444);
  ND2 NAND2_897(g11994,g8310,g8365);
  ND2 NAND2_898(g15723,g10775,g13104);
  ND3 NAND3_136(g23978,g572,g21389,g12323);
  ND4 NAND4_142(g13967,g3929,g11225,g3983,g11419);
  ND2 NAND2_899(I12345,g3106,I12344);
  ND2 NAND2_900(I14790,g6167,I14788);
  ND2 NAND2_901(I14516,g10147,g661);
  ND2 NAND2_902(g23590,g20682,g11111);
  ND2 NAND2_903(I12849,g4281,I12848);
  ND2 NAND2_904(g12008,g9932,g5798);
  ND4 NAND4_143(g17814,g5579,g14522,g5673,g12563);
  ND2 NAND2_905(g22638,g18957,g2886);
  ND2 NAND2_906(I12848,g4281,g4277);
  ND2 NAND2_907(g12476,g7498,g6704);
  ND3 NAND3_137(g13459,g7479,g11294,g11846);
  ND4 NAND4_144(g21384,g17734,g14686,g17675,g14663);
  ND2 NAND2_908(I23587,g4332,I23585);
  ND2 NAND2_909(g8889,g3684,g4871);
  ND2 NAND2_910(g14038,g11514,g11435);
  ND2 NAND2_911(g23067,g20887,g10721);
  ND2 NAND2_912(g10601,g896,g7397);
  ND4 NAND4_145(g13918,g3259,g11217,g3267,g11350);
  ND4 NAND4_146(g16925,g3574,g13799,g3668,g11576);
  ND2 NAND2_913(g14601,g12318,g6466);
  ND2 NAND2_914(I18538,g14642,I18536);
  ND2 NAND2_915(g8871,I12841,I12842);
  ND2 NAND2_916(I15079,g9827,I15078);
  ND2 NAND2_917(g14677,I16779,I16780);
  ND2 NAND2_918(I12263,g1448,I12261);
  ND2 NAND2_919(g11545,I14498,I14499);
  ND3 NAND3_138(g11444,g6905,g6918,g8733);
  ND2 NAND2_920(g13079,g1312,g11336);
  ND2 NAND2_921(I15078,g9827,g1968);
  ND2 NAND2_922(g12239,I15106,I15107);
  ND2 NAND2_923(g20201,I20468,I20469);
  ND2 NAND2_924(g8500,g3431,g3423);
  ND2 NAND2_925(g14937,g12667,g10421);
  ND2 NAND2_926(g26025,g22405,g24631);
  ND4 NAND4_147(g13086,g6235,g12101,g6346,g10003);
  ND2 NAND2_927(g16681,I17884,I17885);
  ND4 NAND4_148(g17578,g5212,g14399,g5283,g12497);
  ND2 NAND2_928(g12941,g7167,g10537);
  ND2 NAND2_929(g19795,g13600,g16275);
  ND2 NAND2_930(g12185,g9905,g799);
  ND4 NAND4_149(g21402,g17757,g14740,g17716,g14674);
  ND2 NAND2_931(g17586,g14638,g14601);
  ND2 NAND2_932(g11977,g8373,g2476);
  ND2 NAND2_933(g13977,g11610,g11729);
  ND2 NAND2_934(I14530,g8840,g8873);
  ND2 NAND2_935(g8737,I12729,I12730);
  ND2 NAND2_936(g15011,g12716,g12632);
  ND2 NAND2_937(g34227,I32203,I32204);
  ND2 NAND2_938(g14015,g11658,g11747);
  ND2 NAND2_939(g11561,I14517,I14518);
  ND2 NAND2_940(g25172,g5052,g23560);
  ND2 NAND2_941(I22872,g12150,I22871);
  ND2 NAND2_942(g25996,g24601,g22838);
  ND4 NAND4_150(g20170,g16741,g13897,g16687,g13866);
  ND2 NAND2_943(g10556,g7971,g8133);
  ND2 NAND2_944(g13823,g11313,g3774);
  ND2 NAND2_945(I13454,g1959,I13452);
  ND2 NAND2_946(I21992,g7670,g19638);
  ND2 NAND2_947(g14223,g9092,g11858);
  ND2 NAND2_948(g17493,g8659,g14367);
  ND2 NAND2_949(g15959,I17405,I17406);
  ND4 NAND4_151(g27577,g25019,g25002,g24988,g25765);
  ND2 NAND2_950(I15364,g10182,I15363);
  ND3 NAND3_139(g12577,g7051,g5990,g6044);
  ND2 NAND2_951(g14110,g11692,g8906);
  ND2 NAND2_952(g9246,g847,g812);
  ND4 NAND4_152(g15742,g5575,g12093,g5637,g14669);
  ND2 NAND2_953(I23586,g22409,I23585);
  ND2 NAND2_954(g9203,g3706,g3752);
  ND4 NAND4_153(g14740,g5913,g12129,g6031,g12614);
  ND2 NAND2_955(I13382,g269,g246);
  ND2 NAND2_956(I15289,g6697,I15287);
  ND2 NAND2_957(g19358,g15723,g1399);
  ND2 NAND2_958(I13519,g2514,I13518);
  ND3 NAND3_140(g16299,g8160,g8112,g13706);
  ND3 NAND3_141(g31003,g27163,g29497,g19644);
  ND2 NAND2_959(g14953,g12646,g12405);
  ND2 NAND2_960(I15288,g10061,I15287);
  ND2 NAND2_961(I13518,g2514,g2518);
  ND2 NAND2_962(g12083,g2217,g8205);
  ND2 NAND2_963(I15308,g2407,I15306);
  ND2 NAND2_964(g11224,I14290,I14291);
  ND2 NAND2_965(g13288,g10946,g1442);
  ND4 NAND4_154(g15730,g6609,g14556,g6711,g10061);
  ND2 NAND2_966(g14800,g7704,g12443);
  ND2 NAND2_967(I24414,g23751,g14382);
  ND2 NAND2_968(g29046,g27779,g9640);
  ND3 NAND3_142(g13495,g1008,g11786,g7972);
  ND2 NAND2_969(I29261,g29485,g12046);
  ND2 NAND2_970(g24809,g19965,g23132);
  ND2 NAND2_971(I22846,g21228,I22844);
  ND2 NAND2_972(g24808,I23986,I23987);
  ND2 NAND2_973(I13729,g4534,g4537);
  ND2 NAND2_974(g10587,g2421,g7456);
  ND2 NAND2_975(g11374,g9536,g1536);
  ND2 NAND2_976(g28391,g27064,g13637);
  ND2 NAND2_977(g12415,g7496,g5976);
  ND2 NAND2_978(g21287,g14616,g17571);
  ND2 NAND2_979(g19506,g4087,g15825);
  ND2 NAND2_980(g10909,g7304,g1116);
  ND3 NAND3_143(g20733,g14406,g17290,g9509);
  ND4 NAND4_155(g21307,g15719,g13067,g15709,g13040);
  ND2 NAND2_981(g15002,g12609,g10312);
  ND2 NAND2_982(I25243,g490,I25242);
  ND2 NAND2_983(g13260,g1116,g10666);
  ND2 NAND2_984(g14908,g7812,g10491);
  ND2 NAND2_985(g10569,g2287,g7418);
  ND2 NAND2_986(I22929,g12223,g21228);
  ND2 NAND2_987(I15195,g6005,I15193);
  ND2 NAND2_988(I17405,g13378,I17404);
  ND2 NAND2_989(I12344,g3106,g3111);
  ND4 NAND4_156(g14569,g3195,g11194,g3329,g8481);
  ND2 NAND2_990(g11489,g9661,g3618);
  ND2 NAND2_991(g10568,g7328,g7374);
  ND2 NAND2_992(g25895,g1259,g24453);
  ND2 NAND2_993(g16316,g9429,g13518);
  ND2 NAND2_994(g11559,I14509,I14510);
  ND2 NAND2_995(g11424,g9662,g4012);
  ND2 NAND2_996(I13566,g2652,I13564);
  ND2 NAND2_997(g23655,I22793,I22794);
  ND2 NAND2_998(I29271,g12050,I29269);
  ND2 NAND2_999(g9883,g5782,g5774);
  ND2 NAND2_1000(g14123,g10685,g10928);
  ND4 NAND4_157(g15737,g13240,g13115,g7903,g13210);
  ND2 NAND2_1001(g14807,g7738,g12453);
  ND3 NAND3_144(g19903,g13707,g16319,g8227);
  ND2 NAND2_1002(g12115,g1926,g8249);
  ND2 NAND2_1003(g14974,g12744,g12622);
  ND4 NAND4_158(g17790,g6311,g14575,g6322,g10003);
  ND3 NAND3_145(g17137,g13727,g13511,g13527);
  ND2 NAND2_1004(I13139,g6154,g6159);
  ND3 NAND3_146(g11544,g8700,g3990,g4045);
  ND4 NAND4_159(g13544,g7972,g10521,g7549,g1008);
  ND2 NAND2_1005(g24570,g22957,g2941);
  ND2 NAND2_1006(g12052,g7387,g2465);
  ND2 NAND2_1007(g14638,g9626,g12361);
  ND2 NAND2_1008(I15042,g9752,I15041);
  ND2 NAND2_1009(I15255,g1848,I15253);
  ND2 NAND2_1010(I13852,g7397,I13850);
  ND2 NAND2_1011(g14841,g12593,g12443);
  ND3 NAND3_147(g25385,g22369,g1783,g8241);
  ND2 NAND2_1012(g24567,g22957,g2917);
  ND2 NAND2_1013(g11189,I14248,I14249);
  ND2 NAND2_1014(g11679,g8836,g802);
  ND2 NAND2_1015(I23600,g22360,g4322);
  ND3 NAND3_148(g29778,g294,g28444,g23204);
  ND4 NAND4_160(g13124,g10666,g7661,g979,g1061);
  ND2 NAND2_1016(g25888,g914,g24439);
  ND2 NAND2_1017(g31971,g30573,g10511);
  ND2 NAND2_1018(g23210,g18957,g2882);
  ND4 NAND4_161(g16696,g13871,g13855,g14682,g12340);
  ND4 NAND4_162(g20185,g16772,g13928,g16723,g13882);
  ND2 NAND2_1019(g10578,g7174,g6058);
  ND3 NAND3_149(g20675,g14377,g17246,g9442);
  ND2 NAND2_1020(g20092,g11373,g17794);
  ND4 NAND4_163(g14014,g3199,g11217,g3298,g11519);
  ND2 NAND2_1021(g11938,g8259,g2208);
  ND2 NAND2_1022(g10586,g7380,g7418);
  ND4 NAND4_164(g13093,g10649,g7661,g979,g1061);
  ND2 NAND2_1023(g8873,I12849,I12850);
  ND2 NAND2_1024(g8632,g1514,g1500);
  ND2 NAND2_1025(g9538,g1792,g1760);
  ND2 NAND2_1026(I20221,g16272,g11170);
  ND2 NAND2_1027(I12240,g1111,g1105);
  ND2 NAND2_1028(g9509,g5770,g5774);
  ND2 NAND2_1029(g23286,g6875,g20887);
  ND2 NAND2_1030(g25426,g12371,g22369);
  ND2 NAND2_1031(g29672,g28376,g13672);
  ND2 NAND2_1032(g17593,I18537,I18538);
  ND2 NAND2_1033(g14116,g11697,g11584);
  ND2 NAND2_1034(I32185,g33665,g33661);
  ND2 NAND2_1035(I14509,g370,I14508);
  ND2 NAND2_1036(g10041,I13565,I13566);
  ND2 NAND2_1037(g14720,g12593,g10266);
  ND2 NAND2_1038(I32518,g34422,I32516);
  ND3 NAND3_150(g16259,g4743,g13908,g12054);
  ND2 NAND2_1039(I14508,g370,g8721);
  ND3 NAND3_151(g16225,g13544,g13528,g13043);
  ND2 NAND2_1040(g14041,g11610,g11473);
  ND2 NAND2_1041(g21187,g14616,g17364);
  ND2 NAND2_1042(I22710,g11915,g21434);
  ND2 NAND2_1043(g12207,g9887,g5794);
  ND2 NAND2_1044(g23975,I23119,I23120);
  ND2 NAND2_1045(g12539,I15341,I15342);
  ND2 NAND2_1046(I24463,g14437,I24461);
  ND4 NAND4_165(g15753,g6239,g14529,g6351,g10003);
  ND2 NAND2_1047(g12538,I15334,I15335);
  ND2 NAND2_1048(I12262,g1454,I12261);
  ND2 NAND2_1049(I13184,g6505,I13182);
  ND2 NAND2_1050(I14213,g9295,I14211);
  ND4 NAND4_166(g15736,g6295,g14575,g6373,g10003);
  ND4 NAND4_167(g17635,g3542,g13730,g3654,g8542);
  ND2 NAND2_1051(g16069,I17447,I17448);
  ND2 NAND2_1052(g13915,g11566,g11473);
  ND2 NAND2_1053(I22945,g9492,I22944);
  ND2 NAND2_1054(g14142,g11715,g8958);
  ND3 NAND3_152(g33925,g33394,g4462,g4467);
  ND4 NAND4_168(g16657,g3554,g13730,g3625,g11576);
  ND2 NAND2_1055(I14205,g8508,I14204);
  ND3 NAND3_153(g15843,g7922,g7503,g13264);
  ND4 NAND4_169(g14517,g3231,g11217,g3321,g8481);
  ND2 NAND2_1056(g24906,g8743,g23088);
  ND2 NAND2_1057(g26714,g9316,g25175);
  ND2 NAND2_1058(g23666,g20875,g11139);
  ND2 NAND2_1059(I26417,g26519,g14247);
  ND4 NAND4_170(g21363,g17708,g14664,g17640,g14598);
  ND2 NAND2_1060(I32439,g34227,g34220);
  ND2 NAND2_1061(g12100,I14956,I14957);
  ND2 NAND2_1062(I17380,g13336,I17379);
  ND2 NAND2_1063(g24566,g22755,g22713);
  ND2 NAND2_1064(g22711,g19581,g7888);
  ND2 NAND2_1065(g14130,g11621,g8906);
  ND2 NAND2_1066(I18682,g14752,I18680);
  ND2 NAND2_1067(g17474,g14547,g14521);
  ND3 NAND3_154(g28516,g10857,g26105,g27155);
  ND2 NAND2_1068(g11419,I14428,I14429);
  ND2 NAND2_1069(g29097,g9700,g27858);
  ND4 NAND4_171(g15709,g5224,g14399,g5327,g9780);
  ND4 NAND4_172(g27882,g21228,g25307,g26424,g26213);
  ND3 NAND3_155(g11155,g4776,g7892,g9030);
  ND2 NAND2_1070(I14350,g8890,g8848);
  ND2 NAND2_1071(g15708,g7340,g13083);
  ND3 NAND3_156(g12414,g7028,g7041,g10165);
  ND2 NAND2_1072(g13822,g8160,g11306);
  ND3 NAND3_157(g13266,g12440,g9920,g9843);
  ND2 NAND2_1073(g25527,g21294,g23462);
  ND2 NAND2_1074(I12098,g1322,I12096);
  ND2 NAND2_1075(g14727,g12604,g12505);
  ND2 NAND2_1076(I12251,g1124,g1129);
  ND2 NAND2_1077(I22717,g11916,g21434);
  ND2 NAND2_1078(g17492,g8655,g14367);
  ND2 NAND2_1079(I17448,g956,I17446);
  ND2 NAND2_1080(I15167,g9904,I15166);
  ND2 NAND2_1081(I15194,g9935,I15193);
  ND2 NAND2_1082(I17404,g13378,g1472);
  ND2 NAND2_1083(I31985,g33648,I31983);
  ND2 NAND2_1084(g21186,g14616,g17363);
  ND2 NAND2_1085(g23685,I22823,I22824);
  ND2 NAND2_1086(g7223,I11878,I11879);
  ND2 NAND2_1087(g14600,g9564,g12311);
  ND4 NAND4_173(g14781,g6259,g12173,g6377,g12672);
  ND2 NAND2_1088(g24576,g22957,g2902);
  ND4 NAND4_174(g13119,g6625,g12211,g6715,g10061);
  ND2 NAND2_1089(g21417,g11677,g17157);
  ND2 NAND2_1090(g11118,I14170,I14171);
  ND2 NAND2_1091(g12114,g8241,g8146);
  ND4 NAND4_175(g13118,g5897,g12067,g6031,g9935);
  ND2 NAND2_1092(g21334,g14616,g17596);
  ND2 NAND2_1093(g24609,g22850,g22650);
  ND2 NAND2_1094(g20200,I20461,I20462);
  ND2 NAND2_1095(I29295,g29495,g12117);
  ND2 NAND2_1096(g22663,I21977,I21978);
  ND3 NAND3_158(g33299,g608,g32296,g12323);
  ND2 NAND2_1097(g23762,I22900,I22901);
  ND2 NAND2_1098(I15053,g2259,I15051);
  ND2 NAND2_1099(I15254,g10078,I15253);
  ND2 NAND2_1100(g27141,I25846,I25847);
  ND2 NAND2_1101(I25909,g24782,I25907);
  ND2 NAND2_1102(g24798,I23962,I23963);
  ND4 NAND4_176(g14422,g3187,g11194,g3298,g8481);
  ND2 NAND2_1103(g24973,g21272,g23462);
  ND4 NAND4_177(g20184,g16770,g13918,g16719,g13896);
  ND2 NAND2_1104(g23909,g7028,g20739);
  ND2 NAND2_1105(I25908,g26256,I25907);
  ND2 NAND2_1106(g22757,g20114,g7891);
  ND2 NAND2_1107(g12332,I15167,I15168);
  ND2 NAND2_1108(g25019,g20055,g23172);
  ND2 NAND2_1109(g25018,g20107,g23154);
  ND2 NAND2_1110(I18633,g2504,g14713);
  ND4 NAND4_178(g14542,g3582,g11238,g3672,g8542);
  ND2 NAND2_1111(g14021,g11697,g8958);
  ND2 NAND2_1112(g24934,g21283,g23462);
  ND2 NAND2_1113(I25242,g490,g24744);
  ND4 NAND4_179(g17757,g5909,g14549,g6005,g12614);
  ND4 NAND4_180(g10726,g7304,g7661,g979,g1061);
  ND2 NAND2_1114(g23747,I22865,I22866);
  ND3 NAND3_159(g10614,g9024,g8977,g8928);
  ND4 NAND4_181(g27833,g21228,g25282,g26424,g26190);
  ND2 NAND2_1115(g12049,g2208,g8150);
  ND2 NAND2_1116(g10905,g1116,g7304);
  ND2 NAND2_1117(I15166,g9904,g9823);
  ND2 NAND2_1118(g14905,g12785,g7142);
  ND2 NAND2_1119(g12048,g7369,g2040);
  ND4 NAND4_182(g20214,g16854,g13993,g16776,g13967);
  ND2 NAND2_1120(g28109,g27051,g25783);
  ND2 NAND2_1121(g12221,I15079,I15080);
  ND4 NAND4_183(g27613,g24942,g24933,g25048,g26871);
  ND2 NAND2_1122(g11892,g7777,g9086);
  ND2 NAND2_1123(g13892,g11653,g11473);
  ND3 NAND3_160(g13476,g7503,g11336,g11869);
  ND4 NAND4_184(g21416,g17775,g14781,g17744,g14706);
  ND2 NAND2_1124(I13141,g6159,I13139);
  ND2 NAND2_1125(I14249,g8091,I14247);
  ND2 NAND2_1126(I17379,g13336,g1129);
  ND2 NAND2_1127(I17925,g1478,I17923);
  ND2 NAND2_1128(I23949,g23162,g13603);
  ND2 NAND2_1129(g14797,g12593,g12405);
  ND3 NAND3_161(g27273,g10504,g26131,g26105);
  ND2 NAND2_1130(I14482,g655,I14480);
  ND4 NAND4_185(g16687,g3255,g13700,g3325,g11519);
  ND2 NAND2_1131(g13712,g8984,g11283);
  ND4 NAND4_186(g17634,g3219,g11217,g3281,g13877);
  ND2 NAND2_1132(g11914,g8187,g1648);
  ND4 NAND4_187(g17872,g6617,g14602,g6711,g12721);
  ND2 NAND2_1133(g12947,g7184,g10561);
  ND2 NAND2_1134(I14248,g1322,I14247);
  ND2 NAND2_1135(I22944,g9492,g19620);
  ND4 NAND4_188(g8728,g3618,g3661,g3632,g3654);
  ND2 NAND2_1136(I14204,g8508,g3821);
  ND2 NAND2_1137(g25300,g22369,g12018);
  ND3 NAND3_162(g27463,g287,g26330,g23204);
  ND4 NAND4_189(g13907,g3941,g11225,g4023,g11631);
  ND2 NAND2_1138(g28381,g27074,g13621);
  ND2 NAND2_1139(g29057,g27800,g9649);
  ND2 NAND2_1140(g12463,g7513,g6322);
  ND2 NAND2_1141(g14136,g11571,g8906);
  ND2 NAND2_1142(g14408,g6069,g11924);
  ND2 NAND2_1143(g12972,g7209,g10578);
  ND2 NAND2_1144(g28174,g1270,g27059);
  ND3 NAND3_163(g28796,g27858,g7418,g7335);
  ND2 NAND2_1145(g31753,I29314,I29315);
  ND2 NAND2_1146(I22793,g11956,I22792);
  ND3 NAND3_164(g16260,g4888,g13910,g12088);
  ND2 NAND2_1147(g7823,I12218,I12219);
  ND3 NAND3_165(g28840,g27858,g7380,g2287);
  ND3 NAND3_166(g11382,g8644,g6895,g8663);
  ND2 NAND2_1148(I15176,g2661,I15174);
  ND2 NAND2_1149(I12203,g1094,g1135);
  ND3 NAND3_167(g19632,g1413,g1542,g16047);
  ND2 NAND2_1150(I24440,g14411,I24438);
  ND2 NAND2_1151(g11675,g8984,g4912);
  ND4 NAND4_190(g13176,g10715,g7675,g1322,g1404);
  ND2 NAND2_1152(g13092,g1061,g10761);
  ND2 NAND2_1153(g26269,I25243,I25244);
  ND3 NAND3_168(g34550,g626,g34359,g12323);
  ND2 NAND2_1154(g11154,I14212,I14213);
  ND2 NAND2_1155(g29737,g28421,g13779);
  ND3 NAND3_169(g28522,g10857,g26131,g27142);
  ND2 NAND2_1156(g8678,g376,g358);
  ND2 NAND2_1157(g17592,I18530,I18531);
  ND3 NAND3_170(g16893,g10685,g13252,g703);
  ND2 NAND2_1158(g10537,g7138,g5366);
  ND2 NAND2_1159(I14331,g225,I14330);
  ND2 NAND2_1160(g8105,g3068,g3072);
  ND2 NAND2_1161(I31984,g33653,I31983);
  ND2 NAND2_1162(g16713,I17924,I17925);
  ND2 NAND2_1163(I20462,g14187,I20460);
  ND2 NAND2_1164(I29255,g12017,I29253);
  ND2 NAND2_1165(I24462,g23796,I24461);
  ND4 NAND4_191(g17820,g5925,g14549,g6019,g12614);
  ND2 NAND2_1166(g31709,I29285,I29286);
  ND4 NAND4_192(g15752,g5921,g12129,g5983,g14701);
  ND2 NAND2_1167(I29270,g29486,I29269);
  ND2 NAND2_1168(g28949,g27903,g14643);
  ND2 NAND2_1169(I13463,g2380,I13462);
  ND2 NAND2_1170(g31708,I29278,I29279);
  ND4 NAND4_193(g17846,g6271,g14575,g6365,g12672);
  ND2 NAND2_1171(g17396,g7345,g14272);
  ND4 NAND4_194(g14750,g6633,g12137,g6715,g12721);
  ND3 NAND3_171(g24584,g22852,g22836,g22715);
  ND2 NAND2_1172(I14212,g9252,I14211);
  ND2 NAND2_1173(g7167,g5360,g5406);
  ND2 NAND2_1174(g10796,g7537,g7523);
  ND2 NAND2_1175(g20107,g11404,g17794);
  ND2 NAND2_1176(g11906,I14713,I14714);
  ND2 NAND2_1177(I12403,g3813,I12401);
  ND2 NAND2_1178(g16093,I17461,I17462);
  ND3 NAND3_172(g12344,g10093,g7041,g10130);
  ND3 NAND3_173(g13083,g4392,g10590,g4434);
  ND2 NAND2_1179(I32441,g34220,I32439);
  ND2 NAND2_1180(g13284,g10695,g1157);
  ND2 NAND2_1181(g7549,g1018,g1030);
  ND2 NAND2_1182(g25341,g22417,g12047);
  ND2 NAND2_1183(g29722,g28410,g13742);
  ND2 NAND2_1184(g25268,g21124,g23692);
  ND4 NAND4_195(g16875,g3223,g13765,g3317,g11519);
  ND2 NAND2_1185(g7598,I12075,I12076);
  ND2 NAND2_1186(I32758,g25779,I32756);
  ND4 NAND4_196(g14663,g5236,g12002,g5290,g12239);
  ND2 NAND2_1187(g24804,g19916,g23105);
  ND3 NAND3_174(g24652,g22712,g22940,g22757);
  ND4 NAND4_197(g13139,g6589,g12137,g6723,g10061);
  ND4 NAND4_198(g15713,g5571,g14425,g5673,g9864);
  ND2 NAND2_1188(I14369,g8481,I14368);
  ND2 NAND2_1189(g34469,I32517,I32518);
  ND2 NAND2_1190(I15333,g10152,g2116);
  ND3 NAND3_175(g19546,g15969,g10841,g10884);
  ND2 NAND2_1191(g8227,g3770,g3774);
  ND2 NAND2_1192(I14368,g8481,g3303);
  ND2 NAND2_1193(g12028,I14884,I14885);
  ND2 NAND2_1194(g15042,g12806,g10491);
  ND2 NAND2_1195(g21253,g6423,g17482);
  ND2 NAND2_1196(I29277,g29488,g12081);
  ND2 NAND2_1197(g23781,I22937,I22938);
  ND2 NAND2_1198(g13963,g11715,g11584);
  ND4 NAND4_199(g17640,g5264,g14399,g5335,g12497);
  ND2 NAND2_1199(I14229,g979,I14228);
  ND4 NAND4_200(g21351,g15729,g13098,g15720,g13069);
  ND2 NAND2_1200(g26666,g9229,g25144);
  ND2 NAND2_1201(I14228,g979,g8055);
  ND2 NAND2_1202(g15030,g12716,g12680);
  ND4 NAND4_201(g27903,g21228,g25316,g26424,g26218);
  ND3 NAND3_176(g13554,g11336,g7582,g1351);
  ND2 NAND2_1203(I17924,g13378,I17923);
  ND3 NAND3_177(g12491,g7285,g4462,g6961);
  ND3 NAND3_178(g28780,g27742,g7308,g1636);
  ND2 NAND2_1204(I22753,g11937,g21434);
  ND2 NAND2_1205(g11312,g8565,g3794);
  ND2 NAND2_1206(g11200,g8592,g3798);
  ND2 NAND2_1207(g25038,g21331,g23363);
  ND3 NAND3_179(g13115,g1008,g11786,g11294);
  ND2 NAND2_1208(I15052,g9759,I15051);
  ND2 NAND2_1209(g14933,g12700,g12571);
  ND2 NAND2_1210(I14925,g5835,I14923);
  ND2 NAND2_1211(g16155,I17495,I17496);
  ND2 NAND2_1212(g17662,I18634,I18635);
  ND3 NAND3_180(g28820,g27742,g1668,g1592);
  ND2 NAND2_1213(I12546,g194,I12544);
  ND2 NAND2_1214(I17461,g13378,I17460);
  ND2 NAND2_1215(g14851,g7738,g12505);
  ND2 NAND2_1216(g27767,I26367,I26368);
  ND2 NAND2_1217(g9775,g4831,g4681);
  ND4 NAND4_202(g20371,g16956,g14088,g16694,g16660);
  ND2 NAND2_1218(g24951,g199,g23088);
  ND2 NAND2_1219(g24972,g19962,g23172);
  ND2 NAND2_1220(g12767,g4467,g6961);
  ND2 NAND2_1221(g13798,g11280,g3423);
  ND2 NAND2_1222(g11973,g8365,g2051);
  ND2 NAND2_1223(g30580,g29335,g19666);
  ND2 NAND2_1224(g29657,g28363,g13634);
  ND4 NAND4_203(g17779,g6637,g14556,g6704,g12471);
  ND2 NAND2_1225(g11674,g8676,g4674);
  ND2 NAND2_1226(g7879,I12262,I12263);
  ND2 NAND2_1227(g23726,g9559,g21140);
  ND2 NAND2_1228(I20203,g16246,g11147);
  ND2 NAND2_1229(g16524,g13822,g13798);
  ND2 NAND2_1230(g26685,g9264,g25160);
  ND2 NAND2_1231(I14429,g4005,I14427);
  ND2 NAND2_1232(g14574,g12256,g6120);
  ND2 NAND2_1233(g12191,I15052,I15053);
  ND4 NAND4_204(g14452,g3538,g11207,g3649,g8542);
  ND2 NAND2_1234(g11934,g8139,g8187);
  ND2 NAND2_1235(g16119,I17475,I17476);
  ND2 NAND2_1236(I14428,g8595,I14427);
  ND2 NAND2_1237(g12521,g7471,g5969);
  ND4 NAND4_205(g17647,g5905,g14497,g5976,g12614);
  ND2 NAND2_1238(I29313,g29501,g12154);
  ND2 NAND2_1239(g8609,g1171,g1157);
  ND2 NAND2_1240(g19450,g11471,g17794);
  ND2 NAND2_1241(I14765,g9808,I14764);
  ND2 NAND2_1242(g11761,I14610,I14611);
  ND2 NAND2_1243(g22651,g20114,g2873);
  ND2 NAND2_1244(I29285,g29489,I29284);
  ND2 NAND2_1245(g14051,g10323,g11527);
  ND2 NAND2_1246(g14072,g11571,g11483);
  ND4 NAND4_206(g16749,g3957,g13772,g4027,g11631);
  ND2 NAND2_1247(g20163,g16663,g13938);
  ND4 NAND4_207(g15782,g6585,g14556,g6697,g10061);
  ND2 NAND2_1248(I29254,g29482,I29253);
  ND2 NAND2_1249(I15214,g1714,I15212);
  ND4 NAND4_208(g14780,g6275,g12101,g6329,g12423);
  ND2 NAND2_1250(g12045,g1783,g8146);
  ND3 NAND3_181(g10820,g9985,g9920,g9843);
  ND4 NAND4_209(g14820,g6307,g12173,g6315,g12423);
  ND4 NAND4_210(g17513,g3247,g13765,g3325,g8481);
  ND3 NAND3_182(g28827,g27837,g7362,g1862);
  ND2 NAND2_1251(g25531,g22763,g2868);
  ND3 NAND3_183(g15853,g14714,g9417,g12337);
  ND2 NAND2_1252(I15241,g10003,g6351);
  ND3 NAND3_184(g12462,g7051,g7064,g10190);
  ND2 NAND2_1253(g13241,g7503,g10544);
  ND2 NAND2_1254(g25186,g5396,g23602);
  ND2 NAND2_1255(g14691,g12695,g12505);
  ND3 NAND3_185(g25953,g22756,g24570,g22688);
  ND2 NAND2_1256(g8803,g128,g4646);
  ND2 NAND2_1257(g9954,g6128,g6120);
  ND2 NAND2_1258(I22792,g11956,g21434);
  ND2 NAND2_1259(I22967,g21228,I22965);
  ND4 NAND4_211(g13100,g6581,g12137,g6692,g10061);
  ND2 NAND2_1260(g23575,I22711,I22712);
  ND2 NAND2_1261(g20173,g16696,g13972);
  ND2 NAND2_1262(g10929,g1099,g7854);
  ND2 NAND2_1263(g31669,I29254,I29255);
  ND3 NAND3_186(g15864,g14833,g12543,g12487);
  ND2 NAND2_1264(g33669,g33378,g862);
  ND2 NAND2_1265(g25334,g21253,g23756);
  ND4 NAND4_212(g17723,g6597,g14556,g6668,g12721);
  ND2 NAND2_1266(g10583,g7475,g862);
  ND3 NAND3_187(g10928,g8181,g8137,g417);
  ND4 NAND4_213(g15748,g13257,g13130,g7922,g13241);
  ND2 NAND2_1267(g21283,g11291,g17157);
  ND2 NAND2_1268(g9912,I13463,I13464);
  ND2 NAND2_1269(I13045,g5120,I13043);
  ND4 NAND4_214(g20134,g17572,g14542,g17495,g14452);
  ND4 NAND4_215(g13515,g12628,g12588,g12524,g12464);
  ND4 NAND4_216(g13882,g3590,g11207,g3672,g11576);
  ND2 NAND2_1270(g24760,I23918,I23919);
  ND2 NAND2_1271(I23961,g23184,g13631);
  ND2 NAND2_1272(g25216,g6088,g23678);
  ND2 NAND2_1273(g14113,g11626,g11537);
  ND2 NAND2_1274(I24385,g14347,I24383);
  ND2 NAND2_1275(g15036,g12780,g12581);
  ND2 NAND2_1276(g19597,g1199,g15995);
  ND2 NAND2_1277(g12629,g7812,g7142);
  ND2 NAND2_1278(I12877,g4200,I12876);
  ND2 NAND2_1279(I13462,g2380,g2384);
  ND2 NAND2_1280(g8847,g4831,g4681);
  ND3 NAND3_188(g12628,g7074,g6336,g6390);
  ND3 NAND3_189(g22850,g1536,g19581,g10699);
  ND2 NAND2_1281(g11441,g9599,g3267);
  ND2 NAND2_1282(I13140,g6154,I13139);
  ND2 NAND2_1283(I22901,g21228,I22899);
  ND3 NAND3_190(g28786,g27837,g7405,g7322);
  ND2 NAND2_1284(g11206,I14276,I14277);
  ND3 NAND3_191(g16238,g4698,g13883,g12054);
  ND2 NAND2_1285(I14499,g8737,I14497);
  ND2 NAND2_1286(g17412,g14520,g14489);
  ND2 NAND2_1287(I18625,g2079,g14712);
  ND2 NAND2_1288(g14768,g12662,g12571);
  ND2 NAND2_1289(g28945,g27854,g8211);
  ND4 NAND4_217(g14803,g5208,g12059,g5308,g12497);
  ND2 NAND2_1290(I14498,g9020,I14497);
  ND3 NAND3_192(g33679,g33394,g10737,g10308);
  ND2 NAND2_1291(g12147,g8302,g8201);
  ND2 NAND2_1292(I12402,g3808,I12401);
  ND2 NAND2_1293(I15107,g5313,I15105);
  ND2 NAND2_1294(I22823,g11978,I22822);
  ND2 NAND2_1295(I14611,g8678,I14609);
  ND2 NAND2_1296(I14924,g9558,I14923);
  ND2 NAND2_1297(g12370,I15213,I15214);
  ND2 NAND2_1298(g25974,g24576,g22837);
  ND4 NAND4_218(g17716,g5957,g14497,g6027,g12614);
  ND2 NAND2_1299(g15008,g12780,g10341);
  ND2 NAND2_1300(I23971,g490,I23969);
  ND2 NAND2_1301(g25293,g21190,g23726);
  ND2 NAND2_1302(g12151,g8316,g8211);
  ND2 NAND2_1303(g19854,I20222,I20223);
  ND4 NAND4_219(g13940,g11426,g8889,g11707,g8829);
  ND2 NAND2_1304(I22966,g12288,I22965);
  ND2 NAND2_1305(g23949,g7074,g21012);
  ND2 NAND2_1306(g28448,g23975,g27377);
  ND2 NAND2_1307(I15263,g10081,I15262);
  ND2 NAND2_1308(g10552,g2153,g7374);
  ND4 NAND4_220(g8751,g3969,g4012,g3983,g4005);
  ND3 NAND3_193(g15907,g14833,g9417,g12487);
  ND2 NAND2_1309(g22681,I21993,I21994);
  ND2 NAND2_1310(g11135,I14186,I14187);
  ND2 NAND2_1311(I14330,g225,g9966);
  ND2 NAND2_1312(g19916,g3029,g16313);
  ND4 NAND4_221(g16728,g13884,g13870,g14089,g11639);
  ND2 NAND2_1313(g12227,g8418,g8330);
  ND2 NAND2_1314(I14764,g9808,g5821);
  ND2 NAND2_1315(g11962,I14789,I14790);
  ND2 NAND2_1316(I29284,g29489,g12085);
  ND2 NAND2_1317(I31973,g33641,I31972);
  ND2 NAND2_1318(I29304,g12121,I29302);
  ND2 NAND2_1319(I18581,g14678,I18579);
  ND2 NAND2_1320(I26051,g13500,I26049);
  ND2 NAND2_1321(I25847,g24799,I25845);
  ND2 NAND2_1322(I26072,g13517,I26070);
  ND2 NAND2_1323(I11825,g4593,I11824);
  ND2 NAND2_1324(I12876,g4200,g4180);
  ND2 NAND2_1325(g14999,g12739,g12824);
  ND3 NAND3_194(g16304,g4765,g13970,g12054);
  ND2 NAND2_1326(g12044,g1657,g8139);
  ND2 NAND2_1327(I15004,g1700,I15002);
  ND4 NAND4_222(g21509,g17820,g14898,g17647,g17608);
  ND4 NAND4_223(g17765,g6649,g14556,g6719,g12721);
  ND2 NAND2_1328(I14259,g3133,I14257);
  ND2 NAND2_1329(I17495,g13378,I17494);
  ND2 NAND2_1330(g27377,g10685,g25930);
  ND4 NAND4_224(g24926,g20172,g20163,g23357,g13995);
  ND2 NAND2_1331(g25275,g22342,g11991);
  ND2 NAND2_1332(g12301,I15148,I15149);
  ND2 NAND2_1333(I14258,g8154,I14257);
  ND2 NAND2_1334(g12120,g2476,g8273);
  ND4 NAND4_225(g27738,g21228,g25243,g26424,g26148);
  ND2 NAND2_1335(I32440,g34227,I32439);
  ND2 NAND2_1336(g25237,g6434,g23711);
  ND2 NAND2_1337(I15106,g9780,I15105);
  ND2 NAND2_1338(g13273,g1459,g10699);
  ND2 NAND2_1339(g19335,g15717,g1056);
  ND2 NAND2_1340(g10961,g1442,g7876);
  ND3 NAND3_195(g29679,g153,g28353,g23042);
  ND4 NAND4_226(g15729,g5949,g14549,g6027,g9935);
  ND2 NAND2_1341(g14505,g12073,g9961);
  ND2 NAND2_1342(I12287,g1484,g1300);
  ND2 NAND2_1343(I14955,g9620,g6181);
  ND2 NAND2_1344(g19965,g3380,g16424);
  ND3 NAND3_196(g11951,g9166,g847,g703);
  ND4 NAND4_227(g15728,g5200,g14399,g5313,g9780);
  ND2 NAND2_1345(g13951,g10295,g11729);
  ND2 NAND2_1346(I12076,g979,I12074);
  ND2 NAND2_1347(g23047,g482,g20000);
  ND2 NAND2_1348(g13795,g11216,g401);
  ND3 NAND3_197(g28896,g27837,g1936,g1862);
  ND2 NAND2_1349(I14171,g3119,I14169);
  ND2 NAND2_1350(g20871,g14434,g17396);
  ND2 NAND2_1351(I22893,g12189,I22892);
  ND2 NAND2_1352(I12269,g1141,g956);
  ND2 NAND2_1353(I13044,g5115,I13043);
  ND4 NAND4_228(g17775,g6255,g14575,g6351,g12672);
  ND2 NAND2_1354(I22865,g12146,I22864);
  ND2 NAND2_1355(g23756,g9621,g21206);
  ND2 NAND2_1356(g14723,g7704,g12772);
  ND2 NAND2_1357(g23780,I22930,I22931);
  ND2 NAND2_1358(g14433,g12035,g9890);
  ND2 NAND2_1359(I24384,g23721,I24383);
  ND4 NAND4_229(g21350,g15751,g15742,g15735,g13108);
  ND2 NAND2_1360(g16312,g13580,g13574);
  ND2 NAND2_1361(g14104,g11514,g8864);
  ND2 NAND2_1362(I25846,g26212,I25845);
  ND2 NAND2_1363(g14343,g11961,g9670);
  ND2 NAND2_1364(g10971,g7867,g7886);
  ND2 NAND2_1365(g28958,g27833,g8249);
  ND2 NAND2_1366(g14971,g12667,g12581);
  ND4 NAND4_230(g16745,g3594,g13730,g3661,g11389);
  ND2 NAND2_1367(g31748,I29303,I29304);
  ND2 NAND2_1368(g26208,g7975,g24751);
  ND4 NAND4_231(g16813,g3614,g13799,g3625,g8542);
  ND2 NAND2_1369(I22938,g21228,I22936);
  ND2 NAND2_1370(g27824,I26394,I26395);
  ND2 NAND2_1371(g13920,g11621,g11483);
  ND2 NAND2_1372(I17460,g13378,g1300);
  ND2 NAND2_1373(g24591,g22833,g22642);
  ND2 NAND2_1374(g24776,g3040,g23052);
  ND2 NAND2_1375(I14817,g9962,I14816);
  ND2 NAND2_1376(g25236,I24415,I24416);
  ND2 NAND2_1377(I15121,g9910,g2102);
  ND2 NAND2_1378(g34422,I32432,I32433);
  ND3 NAND3_198(g28857,g27779,g1802,g1728);
  ND2 NAND2_1379(g14133,g11692,g11747);
  ND2 NAND2_1380(I12279,g1472,I12277);
  ND2 NAND2_1381(I14532,g8873,I14530);
  ND2 NAND2_1382(g13121,g11117,g8411);
  ND3 NAND3_199(g28793,g27800,g7328,g2153);
  ND2 NAND2_1383(I13403,g2250,I13401);
  ND2 NAND2_1384(I12278,g1467,I12277);
  ND2 NAND2_1385(g24950,g19442,g23154);
  ND2 NAND2_1386(I12469,g405,I12468);
  ND3 NAND3_200(g27931,g25425,g25381,g25780);
  ND3 NAND3_201(g28765,g27800,g7374,g7280);
  ND2 NAND2_1387(g7611,g4057,g4064);
  ND2 NAND2_1388(g14011,g10295,g11473);
  ND4 NAND4_232(g20151,g17598,g14570,g17514,g14519);
  ND2 NAND2_1389(g20172,g16876,g8131);
  ND2 NAND2_1390(I12468,g405,g392);
  ND2 NAND2_1391(g13291,g10715,g1500);
  ND3 NAND3_202(g11173,g4966,g7898,g9064);
  ND2 NAND2_1392(g12190,g8365,g8255);
  ND2 NAND2_1393(g22753,g1536,g19632);
  ND3 NAND3_203(g28504,g758,g27528,g11679);
  ND4 NAND4_233(g21357,g15736,g13109,g15726,g13086);
  ND3 NAND3_204(g31009,g27187,g29503,g19644);
  ND2 NAND2_1394(g14627,g12553,g12772);
  ND2 NAND2_1395(g23357,g20201,g11231);
  ND2 NAND2_1396(g14959,g12695,g12798);
  ND2 NAND2_1397(g14379,g5723,g11907);
  ND2 NAND2_1398(g22650,g7888,g19581);
  ND3 NAND3_205(g11134,g8138,g8240,g8301);
  ND2 NAND2_1399(g23105,g8097,g19887);
  ND2 NAND2_1400(g13134,g11134,g8470);
  ND2 NAND2_1401(g14378,g11979,g9731);
  ND2 NAND2_1402(g7209,g6052,g6098);
  ND2 NAND2_1403(g12024,g8381,g8418);
  ND4 NAND4_234(g17650,g6299,g12101,g6315,g14745);
  ND2 NAND2_1404(g10603,g10077,g9751);
  ND4 NAND4_235(g17736,g5563,g14522,g5659,g12563);
  ND4 NAND4_236(g15798,g6629,g14602,g6704,g14786);
  ND2 NAND2_1405(g25021,g21417,g23363);
  ND2 NAND2_1406(I11824,g4593,g4601);
  ND2 NAND2_1407(g15674,g921,g13110);
  ND2 NAND2_1408(g9310,I13078,I13079);
  ND2 NAND2_1409(I14289,g8282,g3835);
  ND3 NAND3_206(g28298,g10533,g26131,g26990);
  ND2 NAND2_1410(g9663,g128,g4646);
  ND4 NAND4_237(g13927,g3578,g11207,g3632,g11389);
  ND2 NAND2_1411(I17494,g13378,g1448);
  ND2 NAND2_1412(g29118,g27886,g9755);
  ND2 NAND2_1413(I12217,g1437,g1478);
  ND4 NAND4_238(g14730,g5615,g12093,g5623,g12301);
  ND2 NAND2_1414(g22709,g1193,g19611);
  ND2 NAND2_1415(I22822,g11978,g21434);
  ND2 NAND2_1416(g13240,g1046,g10521);
  ND2 NAND2_1417(g24957,g21359,g23462);
  ND2 NAND2_1418(g11491,g9982,g4000);
  ND2 NAND2_1419(g12644,g10233,g4531);
  ND2 NAND2_1420(g11903,g9099,g3712);
  ND2 NAND2_1421(I14816,g9962,g6513);
  ND2 NAND2_1422(I32203,g33937,I32202);
  ND2 NAND2_1423(g23890,g7004,g20682);
  ND3 NAND3_207(g12969,g4388,g7178,g10476);
  ND2 NAND2_1424(I13520,g2518,I13518);
  ND2 NAND2_1425(g20645,g14344,g17243);
  ND2 NAND2_1426(g28856,g27738,g8093);
  ND2 NAND2_1427(g14548,g12208,g5774);
  ND2 NAND2_1428(g17225,g8612,g14367);
  ND4 NAND4_239(g17708,g5216,g14490,g5313,g12497);
  ND2 NAND2_1429(g12197,g7296,g5290);
  ND2 NAND2_1430(g8434,g3080,g3072);
  ND3 NAND3_208(g28512,g10857,g27155,g27142);
  ND2 NAND2_1431(g23552,I22684,I22685);
  ND2 NAND2_1432(g15005,g12667,g12622);
  ND2 NAND2_1433(g14317,g5033,g11862);
  ND2 NAND2_1434(g12411,g7393,g5276);
  ND3 NAND3_209(g8347,g4358,g4349,g4340);
  ND2 NAND2_1435(I15262,g10081,g2273);
  ND2 NAND2_1436(g23778,I22922,I22923);
  ND2 NAND2_1437(g11395,g9601,g3983);
  ND2 NAND2_1438(I13497,g255,g232);
  ND2 NAND2_1439(g11990,g9166,g703);
  ND2 NAND2_1440(g13990,g11669,g11584);
  ND2 NAND2_1441(g23786,I22945,I22946);
  ND2 NAND2_1442(I18487,g14611,I18485);
  ND2 NAND2_1443(g13898,g11621,g11747);
  ND2 NAND2_1444(I22864,g12146,g21228);
  ND4 NAND4_240(g21356,g15780,g15752,g15743,g13118);
  ND2 NAND2_1445(I12373,g3457,I12372);
  ND4 NAND4_241(g14626,g12232,g9852,g12159,g9715);
  ND3 NAND3_210(g24661,g23210,g23195,g22984);
  ND3 NAND3_211(g24547,g22638,g22643,g22754);
  ND2 NAND2_1446(I31972,g33641,g33631);
  ND2 NAND2_1447(g12450,g7738,g10281);
  ND3 NAND3_212(g10775,g7960,g7943,g8470);
  ND2 NAND2_1448(g9295,I13066,I13067);
  ND2 NAND2_1449(g12819,g9848,g6961);
  ND2 NAND2_1450(g12910,g11002,g10601);
  ND3 NAND3_213(g34174,g617,g33851,g12323);
  ND4 NAND4_242(g17792,g6601,g14602,g6697,g12721);
  ND2 NAND2_1451(I22900,g12193,I22899);
  ND2 NAND2_1452(g10737,g6961,g9848);
  ND2 NAND2_1453(g25537,g22763,g2873);
  ND2 NAND2_1454(g12111,g847,g9166);
  ND3 NAND3_214(g28271,g10533,g27004,g26990);
  ND2 NAND2_1455(g13861,g1459,g10671);
  ND2 NAND2_1456(g21331,g11402,g17157);
  ND4 NAND4_243(g13573,g8002,g10544,g7582,g1351);
  ND2 NAND2_1457(g23932,g7051,g20875);
  ND2 NAND2_1458(I14713,g9671,I14712);
  ND3 NAND3_215(g12590,g7097,g7110,g10229);
  ND2 NAND2_1459(g33083,g7805,g32118);
  ND2 NAND2_1460(g11389,I14399,I14400);
  ND2 NAND2_1461(g25492,g12479,g22457);
  ND2 NAND2_1462(g14697,g12662,g12824);
  ND2 NAND2_1463(g9966,I13498,I13499);
  ND2 NAND2_1464(g7184,g5706,g5752);
  ND2 NAND2_1465(g9705,g2619,g2587);
  ND2 NAND2_1466(I14610,g8993,I14609);
  ND2 NAND2_1467(I26368,g14211,I26366);
  ND2 NAND2_1468(I29263,g12046,I29261);
  ND2 NAND2_1469(g11534,g7121,g8958);
  ND2 NAND2_1470(I23602,g4322,I23600);
  ND2 NAND2_1471(g20784,g14616,g17595);
  ND3 NAND3_216(g28736,g27742,g7308,g7252);
  ND4 NAND4_244(g19265,g15721,g15715,g13091,g15710);
  ND4 NAND4_245(g13098,g5933,g12129,g6023,g9935);
  ND2 NAND2_1472(I20487,g16696,I20486);
  ND2 NAND2_1473(g11251,g8438,g3092);
  ND2 NAND2_1474(g25381,g538,g23088);
  ND2 NAND2_1475(I23970,g22202,I23969);
  ND4 NAND4_246(g13462,g12449,g12412,g12342,g12294);
  ND3 NAND3_217(g28843,g27907,g7456,g7387);
  ND3 NAND3_218(g19510,g15969,g10841,g10899);
  ND2 NAND2_1476(g20181,g13252,g16846);
  ND2 NAND2_1477(g12019,g7322,g1906);
  ND4 NAND4_247(g17598,g3949,g13824,g4027,g8595);
  ND2 NAND2_1478(g12196,g8764,g4688);
  ND2 NAND2_1479(g11997,g2319,g8316);
  ND2 NAND2_1480(I20469,g16728,I20467);
  ND2 NAND2_1481(I21994,g19638,I21992);
  ND2 NAND2_1482(I12242,g1105,I12240);
  ND3 NAND3_219(g12526,g10194,g7110,g10213);
  ND4 NAND4_248(g15725,g5603,g14522,g5681,g9864);
  ND2 NAND2_1483(I20468,g16663,I20467);
  ND2 NAND2_1484(g29154,g27937,g9835);
  ND4 NAND4_249(g21433,g17792,g14830,g17765,g14750);
  ND2 NAND2_1485(I22892,g12189,g21228);
  ND2 NAND2_1486(g19442,g11431,g17794);
  ND2 NAND2_1487(g12402,g7704,g10266);
  ND2 NAND2_1488(g10611,g10115,g9831);
  ND2 NAND2_1489(I13111,g5813,I13109);
  ND2 NAND2_1490(g13871,g4955,g11834);
  ND2 NAND2_1491(I23919,g9333,I23917);
  ND2 NAND2_1492(I18486,g1677,I18485);
  ND3 NAND3_220(g28259,g10504,g26987,g26973);
  ND2 NAND2_1493(g14924,g12558,g12505);
  ND2 NAND2_1494(I22712,g21434,I22710);
  ND2 NAND2_1495(g17656,I18626,I18627);
  ND2 NAND2_1496(I20187,g16272,g1333);
  ND4 NAND4_250(g15744,g6641,g14602,g6719,g10061);
  ND2 NAND2_1497(I17476,g1105,I17474);
  ND2 NAND2_1498(I23918,g23975,I23917);
  ND2 NAND2_1499(I18580,g1945,I18579);
  ND2 NAND2_1500(I26050,g25997,I26049);
  ND2 NAND2_1501(I13384,g246,I13382);
  ND2 NAND2_1502(g12001,I14854,I14855);
  ND2 NAND2_1503(I13067,g4304,I13065);
  ND2 NAND2_1504(I12841,g4222,I12840);
  ND2 NAND2_1505(I11877,g4388,g4430);
  ND2 NAND2_1506(g10529,g1592,g7308);
  ND2 NAND2_1507(g13628,g3372,g11107);
  ND2 NAND2_1508(g23850,g12185,g19462);
  ND2 NAND2_1509(g13911,g11834,g4917);
  ND2 NAND2_1510(I18531,g14640,I18529);
  ND2 NAND2_1511(g17364,g8639,g14367);
  ND3 NAND3_221(g28955,g27837,g1936,g7362);
  ND2 NAND2_1512(I14277,g3484,I14275);
  ND2 NAND2_1513(I21977,g7680,I21976);
  ND4 NAND4_251(g14696,g5567,g12093,g5685,g12563);
  ND2 NAND2_1514(I24363,g23687,g14320);
  ND2 NAND2_1515(g8163,g3419,g3423);
  ND3 NAND3_222(g15962,g14833,g9417,g9340);
  ND2 NAND2_1516(g14764,g7738,g12798);
  ND2 NAND2_1517(g11591,I14531,I14532);
  ND3 NAND3_223(g21011,g14504,g17399,g9629);
  ND2 NAND2_1518(I15147,g9864,g5659);
  ND2 NAND2_1519(g12066,I14924,I14925);
  ND2 NAND2_1520(I20486,g16696,g16757);
  ND2 NAND2_1521(g24943,g20068,g23172);
  ND3 NAND3_224(g20644,g14342,g17220,g9372);
  ND2 NAND2_1522(g27876,I26418,I26419);
  ND3 NAND3_225(g15833,g14714,g12378,g12337);
  ND2 NAND2_1523(I13402,g2246,I13401);
  ND2 NAND2_1524(g11355,g9551,g3310);
  ND3 NAND3_226(g28994,g27907,g2495,g7424);
  ND2 NAND2_1525(g14868,g12755,g12680);
  ND2 NAND2_1526(g17571,g8579,g14367);
  ND2 NAND2_1527(I11866,g4401,I11864);
  ND4 NAND4_252(g27854,g21228,g25283,g26424,g26195);
  ND2 NAND2_1528(g25062,g21403,g23363);
  ND2 NAND2_1529(I20223,g11170,I20221);
  ND2 NAND2_1530(g16507,g13797,g13764);
  ND2 NAND2_1531(g11858,g9014,g3010);
  ND2 NAND2_1532(I14352,g8848,I14350);
  ND2 NAND2_1533(I17883,g13336,g1135);
  ND2 NAND2_1534(g11172,g8478,g3096);
  ND3 NAND3_227(g12511,g7028,g5644,g5698);
  ND2 NAND2_1535(g22687,g19560,g7870);
  ND2 NAND2_1536(g7885,I12270,I12271);
  ND2 NAND2_1537(g11996,g7280,g2197);
  ND4 NAND4_253(g17495,g3566,g13730,g3668,g8542);
  ND2 NAND2_1538(g23379,g20216,g11248);
  ND2 NAND2_1539(I14170,g8389,I14169);
  ND2 NAND2_1540(I13077,g5462,g5467);
  ND2 NAND2_1541(g23112,g21024,g10733);
  ND3 NAND3_228(g20870,g14432,g17315,g9567);
  ND4 NAND4_254(g17816,g6657,g14602,g6668,g10061);
  ND2 NAND2_1542(g14258,g9203,g11903);
  ND2 NAND2_1543(g11394,g9600,g3661);
  ND2 NAND2_1544(g22643,g20136,g18954);
  ND2 NAND2_1545(g34051,I31973,I31974);
  ND4 NAND4_255(g21386,g15798,g15788,g15782,g13139);
  ND2 NAND2_1546(I18587,g2370,g14679);
  ND4 NAND4_256(g21603,g17872,g14987,g17723,g17689);
  ND2 NAND2_1547(I14853,g9433,g5142);
  ND2 NAND2_1548(g27550,g24943,g25772);
  ND2 NAND2_1549(g9485,g1657,g1624);
  ND2 NAND2_1550(g14069,g11653,g8864);
  ND2 NAND2_1551(g22668,g20219,g2912);
  ND2 NAND2_1552(g10602,g7411,g7451);
  ND3 NAND3_229(g11446,g8700,g6941,g8734);
  ND2 NAND2_1553(g14810,g12700,g10312);
  ND2 NAND2_1554(g15033,g12806,g7142);
  ND2 NAND2_1555(g12287,g8381,g2587);
  ND4 NAND4_257(g21429,g17788,g14803,g17578,g17520);
  ND4 NAND4_258(g17669,g3570,g11238,g3632,g13902);
  ND2 NAND2_1556(g12307,g7395,g5983);
  ND2 NAND2_1557(g14879,g12646,g10266);
  ND2 NAND2_1558(I13066,g4308,I13065);
  ND4 NAND4_259(g17668,g3235,g13765,g3310,g13877);
  ND2 NAND2_1559(g23428,g13945,g20522);
  ND2 NAND2_1560(g13058,g10544,g1312);
  ND3 NAND3_230(g28977,g27937,g2629,g2555);
  ND2 NAND2_1561(g12431,I15254,I15255);
  ND2 NAND2_1562(g20979,g5385,g17309);
  ND3 NAND3_231(g28783,g27779,g7315,g1728);
  ND2 NAND2_1563(g20055,g11269,g17794);
  ND4 NAND4_260(g20111,g17513,g14517,g17468,g14422);
  ND2 NAND2_1564(g17525,g14600,g14574);
  ND2 NAND2_1565(I13511,g2093,I13509);
  ND2 NAND2_1566(g12341,g7512,g5308);
  ND2 NAND2_1567(g28823,g27738,g14565);
  ND2 NAND2_1568(I14276,g8218,I14275);
  ND2 NAND2_1569(I21976,g7680,g19620);
  ND2 NAND2_1570(g16291,g13551,g13545);
  ND2 NAND2_1571(I23985,g22182,g482);
  ND2 NAND2_1572(g13281,g10916,g1099);
  ND2 NAND2_1573(g27670,g25172,g26666);
  ND2 NAND2_1574(g22713,g20114,g2890);
  ND2 NAND2_1575(g11957,g8205,g8259);
  ND4 NAND4_261(g28336,g27064,g24756,g27163,g19644);
  ND2 NAND2_1576(I32202,g33937,g33670);
  ND2 NAND2_1577(g13739,g11773,g11261);
  ND3 NAND3_232(g25396,g22384,g2208,g8259);
  ND3 NAND3_233(g28966,g27858,g2361,g7380);
  ND2 NAND2_1578(g14918,g12646,g12772);
  ND4 NAND4_262(g20150,g17705,g17669,g17635,g14590);
  ND2 NAND2_1579(g14079,g11626,g11763);
  ND4 NAND4_263(g17705,g3586,g13799,g3661,g13902);
  ND2 NAND2_1580(g8292,g218,g215);
  ND2 NAND2_1581(g14599,g12207,g9739);
  ND2 NAND2_1582(I12253,g1129,I12251);
  ND4 NAND4_264(g17679,g5611,g14425,g5681,g12563);
  ND2 NAND2_1583(g7869,I12252,I12253);
  ND2 NAND2_1584(g10598,g7191,g6404);
  ND4 NAND4_265(g15788,g6613,g12211,g6675,g14786);
  ND2 NAND2_1585(I18579,g1945,g14678);
  ND4 NAND4_266(g14598,g5248,g12002,g5331,g12497);
  ND2 NAND2_1586(I14733,g9732,g5475);
  ND2 NAND2_1587(g15829,g4112,g13831);
  ND4 NAND4_267(g17686,g6251,g14529,g6322,g12672);
  ND2 NAND2_1588(I12372,g3457,g3462);
  ND2 NAND2_1589(g14817,g12711,g12622);
  ND3 NAND3_234(g28288,g10533,g26105,g27004);
  ND2 NAND2_1590(g19913,g11430,g17794);
  ND2 NAND2_1591(g19614,g1542,g16047);
  ND2 NAND2_1592(g22875,g20516,g2980);
  ND2 NAND2_1593(g25020,g21377,g23462);
  ND2 NAND2_1594(g7442,g896,g890);
  ND2 NAND2_1595(g24917,g19913,g23172);
  ND2 NAND2_1596(g10561,g7157,g5712);
  ND4 NAND4_268(g27468,g24951,g24932,g24925,g26852);
  ND2 NAND2_1597(I22921,g14677,g21284);
  ND2 NAND2_1598(g27306,g24787,g26235);
  ND2 NAND2_1599(g19530,g15829,g10841);
  ND2 NAND2_1600(g12286,I15129,I15130);
  ND2 NAND2_1601(g14656,g12553,g12405);
  ND2 NAND2_1602(g9177,g3355,g3401);
  ND2 NAND2_1603(g22837,g20219,g2907);
  ND2 NAND2_1604(g12306,g7394,g5666);
  ND2 NAND2_1605(I26461,g14306,I26459);
  ND2 NAND2_1606(I24416,g14382,I24414);
  ND4 NAND4_269(g16604,g3251,g11194,g3267,g13877);
  ND2 NAND2_1607(I22799,g11960,g21434);
  ND4 NAND4_270(g13551,g11812,g7479,g7903,g10521);
  ND2 NAND2_1608(g10336,I13750,I13751);
  ND2 NAND2_1609(g28976,g27903,g8273);
  ND2 NAND2_1610(I14712,g9671,g5128);
  ND2 NAND2_1611(I13335,g1687,I13334);
  ND4 NAND4_271(g16770,g3263,g13765,g3274,g8481);
  ND2 NAND2_1612(g8561,g3782,g3774);
  ND2 NAND2_1613(I22973,g9657,I22972);
  ND2 NAND2_1614(g26248,I25220,I25221);
  ND2 NAND2_1615(g12187,I15042,I15043);
  ND2 NAND2_1616(I29262,g29485,I29261);
  ND3 NAND3_235(g11490,g8666,g3639,g3694);
  ND2 NAND2_1617(I26393,g26488,g14227);
  NR2 NOR2_0(g30249,g5297,g28982);
  NR2 NOR2_1(g33141,g32099,g8400);
  NR2 NOR2_2(g13824,g8623,g11702);
  NR2 NOR2_3(g27479,g9056,g26616);
  NR2 NOR2_4(g12479,g2028,g8310);
  NR2 NOR2_5(g20854,g5381,g17243);
  NR2 NOR2_6(g33135,g32090,g8350);
  NR4 NOR4_0(g7675,g1554,g1559,g1564,g1548);
  NR4 NOR4_1(g12486,g9055,g9013,g8957,g8905);
  NR2 NOR2_7(g9694,g1936,g1862);
  NR2 NOR2_8(g8906,g3530,g3522);
  NR2 NOR2_9(g14816,g10166,g12252);
  NR2 NOR2_10(g12223,g2051,g8365);
  NR2 NOR2_11(g14687,g5352,g12166);
  NR2 NOR2_12(g14752,g12540,g10040);
  NR2 NOR2_13(g16272,g13580,g11189);
  NR2 NOR2_14(g22524,g19720,g1361);
  NR2 NOR2_15(g25778,g25459,g25420);
  NR2 NOR2_16(g26212,g23837,g25408);
  NR2 NOR2_17(g17194,g11039,g13480);
  NR2 NOR2_18(g14392,g12114,g9537);
  NR2 NOR2_19(g13700,g3288,g11615);
  NR2 NOR2_20(g11658,g8021,g3506);
  NR2 NOR2_21(g15718,g13858,g11330);
  NR3 NOR3_0(g10488,g4616,g7133,g10336);
  NR3 NOR3_1(g29107,g6203,g7791,g26977);
  NR3 NOR3_2(g10893,g1189,g7715,g7749);
  NR2 NOR2_22(g25932,g7680,g24528);
  NR2 NOR2_23(g29141,g9374,g27999);
  NR2 NOR2_24(g14713,g12483,g9974);
  NR2 NOR2_25(g31507,g9064,g29556);
  NR2 NOR2_26(g15099,g13191,g12869);
  NR2 NOR2_27(g11527,g8165,g8114);
  NR3 NOR3_3(g32715,g31327,I30261,I30262);
  NR2 NOR2_28(g15098,g13191,g6927);
  NR2 NOR2_29(g30148,g28799,g7335);
  NR2 NOR2_30(g23602,g9672,g20979);
  NR2 NOR2_31(g28470,g8021,g27617);
  NR2 NOR2_32(g16220,g13499,g4939);
  NR2 NOR2_33(g14679,g12437,g9911);
  NR2 NOR2_34(g23955,g2823,g18890);
  NR2 NOR2_35(g33163,g32099,g7809);
  NR2 NOR2_36(g24619,g23554,g23581);
  NR2 NOR2_37(g14188,g9162,g12259);
  NR2 NOR2_38(g14124,g8830,g11083);
  NR2 NOR2_39(g14678,g12432,g9907);
  NR2 NOR2_40(g16246,g13551,g11169);
  NR2 NOR2_41(g12117,g10113,g9755);
  NR2 NOR2_42(g29361,g7553,g28174);
  NR2 NOR2_43(g15140,g12887,g13680);
  NR2 NOR2_44(g14093,g8833,g11083);
  NR2 NOR2_45(g15061,g6815,g13394);
  NR3 NOR3_4(g13910,g4899,g4975,g11173);
  NR2 NOR2_46(g13202,g8347,g10511);
  NR2 NOR2_47(g12123,g6856,g2748);
  NR2 NOR2_48(g27772,g7297,g25839);
  NR2 NOR2_49(g12772,g5188,g9300);
  NR2 NOR2_50(g31121,g4776,g29540);
  NR2 NOR2_51(g23918,g2799,g21382);
  NR2 NOR2_52(g15162,g13809,g12904);
  NR2 NOR2_53(g11384,g8538,g8540);
  NR2 NOR2_54(g23079,g8390,g19965);
  NR2 NOR2_55(g29106,g9451,g28020);
  NR2 NOR2_56(g13094,g7487,g10762);
  NR2 NOR2_57(g26603,g24908,g24900);
  NR3 NOR3_5(g29033,g5511,g7738,g28010);
  NR2 NOR2_58(g15628,g11907,g14228);
  NR3 NOR3_6(g32520,g31554,I30054,I30055);
  NR2 NOR2_59(g17239,g11119,g13518);
  NR3 NOR3_7(g31134,g8033,g29679,g24732);
  NR2 NOR2_60(g33134,g7686,g32057);
  NR2 NOR2_61(g16227,g1554,g13574);
  NR2 NOR2_62(g27007,g5706,g25821);
  NR2 NOR2_63(g31506,g4793,g29540);
  NR2 NOR2_64(g15071,g6831,g13416);
  NR2 NOR2_65(g15147,g13716,g12892);
  NR3 NOR3_8(g15754,g341,g7440,g13385);
  NR2 NOR2_66(g14037,g8748,g11083);
  NR2 NOR2_67(g15825,g7666,g13217);
  NR2 NOR2_68(g16044,g10961,g13861);
  NR2 NOR2_69(g27720,g9253,g25791);
  NR2 NOR2_70(g14419,g12152,g9546);
  NR2 NOR2_71(g29012,g5863,g28020);
  NR2 NOR2_72(g15151,g13745,g7027);
  NR2 NOR2_73(g14418,g12151,g9594);
  NR2 NOR2_74(g10266,g5188,g5180);
  NR2 NOR2_75(g25958,g7779,g24609);
  NR3 NOR3_9(g32296,g9044,g31509,g12259);
  NR2 NOR2_76(g31491,g8938,g29725);
  NR2 NOR2_77(g11280,g8647,g3408);
  NR2 NOR2_78(g25944,g7716,g24591);
  NR2 NOR2_79(g29359,g7528,g28167);
  NR2 NOR2_80(g12806,g9472,g9407);
  NR2 NOR2_81(g14194,g5029,g10515);
  NR2 NOR2_82(g19413,g17151,g14221);
  NR3 NOR3_10(g24953,g10262,g23978,g12259);
  NR2 NOR2_83(g15059,g12839,g13350);
  NR2 NOR2_84(g26298,g8297,g24825);
  NR2 NOR2_85(g30129,g28739,g14537);
  NR2 NOR2_86(g15058,g12838,g13350);
  NR3 NOR3_11(g11231,g7928,g4801,g4793);
  NR2 NOR2_87(g17284,g9253,g14317);
  NR2 NOR2_88(g12193,g2342,g8316);
  NR2 NOR2_89(g11885,g7153,g7167);
  NR3 NOR3_12(g29173,g9259,g27999,g7704);
  NR2 NOR2_90(g14313,g12016,g9250);
  NR2 NOR2_91(g28476,g27627,g26547);
  NR2 NOR2_92(g16226,g8052,g13545);
  NR2 NOR2_93(g11763,g3881,g8172);
  NR2 NOR2_94(g25504,g22550,g7222);
  NR2 NOR2_95(g15120,g12873,g13605);
  NR3 NOR3_13(g32910,g31327,I30468,I30469);
  NR2 NOR2_96(g25317,g9766,g23782);
  NR2 NOR2_97(g10808,g8509,g7611);
  NR2 NOR2_98(g15146,g13716,g7003);
  NR2 NOR2_99(g14036,g8725,g11083);
  NR2 NOR2_100(g34737,g34706,g30003);
  NR2 NOR2_101(g12437,g2319,g8267);
  NR2 NOR2_102(g27703,g9607,g25791);
  NR2 NOR2_103(g20000,g13661,g16264);
  NR2 NOR2_104(g13480,g3017,g11858);
  NR2 NOR2_105(g14642,g12374,g9829);
  NR2 NOR2_106(g12347,g9321,g9274);
  NR2 NOR2_107(g14064,g9214,g12259);
  NR2 NOR2_108(g13076,g7443,g10741);
  NR2 NOR2_109(g33098,g31997,g4616);
  NR3 NOR3_14(g28519,g8011,g27602,g10295);
  NR4 NOR4_2(g12821,g7132,g10223,g7149,g10261);
  NR2 NOR2_110(g27063,g26485,g26516);
  NR2 NOR2_111(g24751,g3034,g23105);
  NR2 NOR2_112(g29903,g6928,g28484);
  NR2 NOR2_113(g11773,g8883,g4785);
  NR2 NOR2_114(g27516,g9180,g26657);
  NR2 NOR2_115(g33140,g7693,g32072);
  NR2 NOR2_116(g13341,g7863,g10762);
  NR2 NOR2_117(g12137,g6682,g7097);
  NR2 NOR2_118(g13670,g8123,g10756);
  NR3 NOR3_15(g10555,g7227,g4601,g4608);
  NR2 NOR2_119(g20841,g17847,g12027);
  NR3 NOR3_16(g23042,g16581,g19462,g10685);
  NR2 NOR2_120(g14712,g12479,g9971);
  NR2 NOR2_121(g13335,g7851,g10741);
  NR2 NOR2_122(g19890,g16987,g8058);
  NR2 NOR2_123(g14914,g12822,g12797);
  NR2 NOR2_124(g24391,g22190,g14645);
  NR2 NOR2_125(g15127,g12879,g13605);
  NR2 NOR2_126(g30271,g7041,g29008);
  NR2 NOR2_127(g23124,g8443,g20011);
  NR2 NOR2_128(g23678,g9809,g21190);
  NR2 NOR2_129(g16024,g14216,g11890);
  NR2 NOR2_130(g12208,g10096,g5759);
  NR2 NOR2_131(g33447,g31978,g7643);
  NR2 NOR2_132(g26330,g8631,g24825);
  NR2 NOR2_133(g23686,g2767,g21066);
  NR2 NOR2_134(g20014,g17096,g11244);
  NR2 NOR2_135(g33162,g4859,g32072);
  NR2 NOR2_136(g29898,g6895,g28458);
  NR2 NOR2_137(g12453,g9444,g5527);
  NR2 NOR2_138(g15095,g13177,g12866);
  NR2 NOR2_139(g29191,g7738,g28010);
  NR2 NOR2_140(g19778,g16268,g1061);
  NR2 NOR2_141(g11618,g8114,g8070);
  NR2 NOR2_142(g14382,g9390,g11139);
  NR2 NOR2_143(g14176,g9044,g12259);
  NR2 NOR2_144(g14092,g8774,g11083);
  NR2 NOR2_145(g19999,g16232,g13742);
  NR2 NOR2_146(g22400,g19345,g15718);
  NR2 NOR2_147(g20720,g17847,g9299);
  NR3 NOR3_17(g11469,g650,g9903,g645);
  NR2 NOR2_148(g12593,g9234,g5164);
  NR2 NOR2_149(g12346,g9931,g9933);
  NR3 NOR3_18(g24720,g1322,g23051,g19793);
  NR2 NOR2_150(g11039,g9056,g9092);
  NR2 NOR2_151(g11306,g3412,g8647);
  NR2 NOR2_152(g30132,g28789,g7362);
  NR2 NOR2_153(g22539,g1030,g19699);
  NR2 NOR2_154(g8958,g3881,g3873);
  NR2 NOR2_155(g33147,g32090,g7788);
  NR2 NOR2_156(g9061,g3401,g3361);
  NR2 NOR2_157(g19932,g3376,g16296);
  NR2 NOR2_158(g25887,g24984,g11706);
  NR2 NOR2_159(g15089,g13144,g12861);
  NR2 NOR2_160(g15088,g13144,g6874);
  NR3 NOR3_19(g13937,g8883,g4785,g11155);
  NR3 NOR3_20(g21277,g9417,g9340,g17467);
  NR2 NOR2_161(g29032,g9300,g27999);
  NR2 NOR2_162(g15126,g12878,g13605);
  NR2 NOR2_163(g11666,g8172,g8125);
  NR2 NOR2_164(g16581,g13756,g8086);
  NR2 NOR2_165(g11363,g8626,g8751);
  NR2 NOR2_166(g11217,g8531,g6875);
  NR2 NOR2_167(g31318,g4785,g29697);
  NR2 NOR2_168(g12711,g6209,g9326);
  NR3 NOR3_21(g8177,g4966,g4991,g4983);
  NR2 NOR2_169(g30171,g28880,g7431);
  NR2 NOR2_170(g17515,g13221,g10828);
  NR2 NOR2_171(g15060,g13350,g6814);
  NR3 NOR3_22(g12492,g7704,g5170,g5164);
  NR2 NOR2_172(g26545,g24881,g24855);
  NR2 NOR2_173(g27982,g7212,g25856);
  NR2 NOR2_174(g27381,g8075,g26657);
  NR2 NOR2_175(g14415,g12147,g9590);
  NR2 NOR2_176(g13110,g7841,g10741);
  NR3 NOR3_23(g26598,g8990,g13756,g24732);
  NR2 NOR2_177(g33146,g4669,g32057);
  NR2 NOR2_178(g29071,g5873,g28020);
  NR2 NOR2_179(g29370,g28585,g28599);
  NR2 NOR2_180(g33427,g10278,g31950);
  NR2 NOR2_181(g22399,g1367,g19720);
  NR2 NOR2_182(g10312,g5881,g5873);
  NR2 NOR2_183(g15055,g6808,g13350);
  NR2 NOR2_184(g15070,g6829,g13416);
  NR2 NOR2_185(g30159,g28799,g14589);
  NR2 NOR2_186(g23560,g9607,g20838);
  NR2 NOR2_187(g12483,g2453,g8324);
  NR2 NOR2_188(g11216,g7998,g8037);
  NR2 NOR2_189(g10799,g347,g7541);
  NR2 NOR2_190(g12553,g5170,g9206);
  NR2 NOR2_191(g23642,g9733,g21124);
  NR2 NOR2_192(g15067,g12842,g13394);
  NR2 NOR2_193(g15094,g13177,g12865);
  NR2 NOR2_194(g30144,g28789,g7322);
  NR2 NOR2_195(g24453,g7446,g22325);
  NR2 NOR2_196(g15150,g12895,g13745);
  NR2 NOR2_197(g31127,g4966,g29556);
  NR3 NOR3_24(g13908,g4709,g8796,g11155);
  NR2 NOR2_198(g12252,g9995,g10185);
  NR2 NOR2_199(g26309,g8575,g24825);
  NR2 NOR2_200(g11747,g3530,g8114);
  NR2 NOR2_201(g13568,g8046,g12527);
  NR2 NOR2_202(g16066,g10929,g13307);
  NR2 NOR2_203(g16231,g13515,g4771);
  NR2 NOR2_204(g33103,g32176,g31212);
  NR2 NOR2_205(g19793,g16292,g1404);
  NR2 NOR2_206(g33095,g31997,g7236);
  NR2 NOR2_207(g12847,g6838,g10430);
  NR2 NOR2_208(g25144,g5046,g23623);
  NR2 NOR2_209(g13772,g3990,g11702);
  NR2 NOR2_210(g28515,g3881,g27635);
  NR2 NOR2_211(g28414,g27467,g26347);
  NR2 NOR2_212(g30288,g7087,g29073);
  NR2 NOR2_213(g26976,g5016,g25791);
  NR2 NOR2_214(g29146,g6565,g26994);
  NR2 NOR2_215(g12851,g6846,g10430);
  NR2 NOR2_216(g14539,g11977,g9833);
  NR2 NOR2_217(g9649,g2227,g2153);
  NR2 NOR2_218(g14538,g11973,g9828);
  NR2 NOR2_219(g28584,g7121,g27635);
  NR2 NOR2_220(g16287,g13622,g11144);
  NR2 NOR2_221(g33089,g31978,g4322);
  NR2 NOR2_222(g15102,g14591,g6954);
  NR2 NOR2_223(g15157,g13782,g12900);
  NR2 NOR2_224(g33088,g31997,g7224);
  NR2 NOR2_225(g22514,g19699,g1018);
  NR2 NOR2_226(g12311,g6109,g10136);
  NR2 NOR2_227(g15066,g12841,g13394);
  NR2 NOR2_228(g24575,g23498,g23514);
  NR2 NOR2_229(g30260,g7018,g28982);
  NR2 NOR2_230(g23883,g2779,g21067);
  NR2 NOR2_231(g26865,g25328,g25290);
  NR2 NOR2_232(g31126,g7928,g29540);
  NR2 NOR2_233(g16268,g7913,g13121);
  NR2 NOR2_234(g12780,g9402,g9326);
  NR2 NOR2_235(g14515,g12225,g9761);
  NR2 NOR2_236(g14414,g12145,g9639);
  NR2 NOR2_237(g11493,g8964,g8967);
  NR2 NOR2_238(g25954,g7750,g24591);
  NR2 NOR2_239(g23729,g17482,g21206);
  NR2 NOR2_240(g20982,g17929,g12065);
  NR2 NOR2_241(g19880,g16201,g13634);
  NR2 NOR2_242(g27731,g9229,g25791);
  NR2 NOR2_243(g12846,g6837,g10430);
  NR2 NOR2_244(g22535,g19699,g1030);
  NR2 NOR2_245(g13806,g11245,g4076);
  NR2 NOR2_246(g29889,g6905,g28471);
  NR2 NOR2_247(g26686,g23678,g25189);
  NR2 NOR2_248(g13517,g8541,g12692);
  NR2 NOR2_249(g20390,g17182,g14257);
  NR2 NOR2_250(g29181,g6573,g26994);
  NR2 NOR2_251(g21284,g16646,g9690);
  NR2 NOR2_252(g26267,g8033,g24732);
  NR2 NOR2_253(g12405,g9374,g5180);
  NR2 NOR2_254(g16210,g13479,g4894);
  NR2 NOR2_255(g15054,g12837,g13350);
  NR2 NOR2_256(g27046,g7544,g25888);
  NR2 NOR2_257(g15156,g13782,g7050);
  NR2 NOR2_258(g30294,g7110,g29110);
  NR2 NOR2_259(g12046,g10036,g9640);
  NR2 NOR2_260(g14399,g5297,g12598);
  NR2 NOR2_261(g11006,g7686,g7836);
  NR2 NOR2_262(g12113,g1648,g8187);
  NR2 NOR2_263(g28106,g7812,g26994);
  NR2 NOR2_264(g25189,g6082,g23726);
  NR2 NOR2_265(g27827,g9456,g25839);
  NR2 NOR2_266(g9586,g1668,g1592);
  NR2 NOR2_267(g19887,g3025,g16275);
  NR2 NOR2_268(g29497,g22763,g28241);
  NR2 NOR2_269(g27769,g9434,g25805);
  NR2 NOR2_270(g15131,g12881,g13638);
  NR2 NOR2_271(g27768,g9264,g25805);
  NR2 NOR2_272(g30160,g28846,g7387);
  NR2 NOR2_273(g33094,g31950,g4639);
  NR2 NOR2_274(g14361,g12079,g9413);
  NR2 NOR2_275(g20183,g17152,g14222);
  NR2 NOR2_276(g28514,g8165,g27617);
  NR2 NOR2_277(g22491,g1361,g19720);
  NR2 NOR2_278(g16479,g14719,g12490);
  NR2 NOR2_279(g27027,g26398,g26484);
  NR2 NOR2_280(g24508,g23577,g23618);
  NR2 NOR2_281(g23052,g8334,g19916);
  NR2 NOR2_282(g12662,g5863,g9274);
  NR2 NOR2_283(g25160,g5390,g23659);
  NR2 NOR2_284(g12249,g5763,g10096);
  NR2 NOR2_285(g11834,g8938,g8822);
  NR2 NOR2_286(g12204,g9927,g10160);
  NR2 NOR2_287(g15143,g6998,g13680);
  NR2 NOR2_288(g30170,g28846,g14615);
  NR2 NOR2_289(g29503,g22763,g28250);
  NR2 NOR2_290(g14033,g8808,g12259);
  NR2 NOR2_291(g12081,g10079,g9694);
  NR2 NOR2_292(g13021,g7544,g10741);
  NR2 NOR2_293(g22521,g1036,g19699);
  NR2 NOR2_294(g27647,g3004,g26616);
  NR2 NOR2_295(g11913,g7197,g9166);
  NR2 NOR2_296(g13913,g8859,g11083);
  NR2 NOR2_297(g27356,g9429,g26657);
  NR2 NOR2_298(g7601,g1322,g1333);
  NR2 NOR2_299(g15168,g13835,g12909);
  NR2 NOR2_300(g27826,g9501,g25821);
  NR2 NOR2_301(g29910,g3990,g28484);
  NR3 NOR3_25(g11607,g8848,g8993,g376);
  NR2 NOR2_302(g14514,g11959,g9760);
  NR2 NOR2_303(g11346,g7980,g7964);
  NR3 NOR3_26(g29070,g5857,g7766,g28020);
  NR2 NOR2_304(g12651,g9269,g5511);
  NR2 NOR2_305(g10421,g6227,g9518);
  NR2 NOR2_306(g30119,g28761,g7315);
  NR2 NOR2_307(g14163,g8997,g12259);
  NR2 NOR2_308(g11797,g8883,g8796);
  NR2 NOR2_309(g19919,g16987,g11205);
  NR2 NOR2_310(g30276,g7074,g29073);
  NR2 NOR2_311(g30285,g7097,g29110);
  NR2 NOR2_312(g19444,g17192,g14295);
  NR2 NOR2_313(g12505,g9444,g9381);
  NR2 NOR2_314(g27717,g9492,g26745);
  NR2 NOR2_315(g9100,g3752,g3712);
  NR2 NOR2_316(g12026,g9417,g9340);
  NR2 NOR2_317(g8984,g4899,g4975);
  NR2 NOR2_318(g14121,g8891,g12259);
  NR2 NOR2_319(g25022,g714,g23324);
  NR2 NOR2_320(g11891,g812,g9166);
  NR2 NOR2_321(g16242,g13529,g4961);
  NR2 NOR2_322(g28491,g8114,g27617);
  NR2 NOR2_323(g33085,g31978,g4311);
  NR2 NOR2_324(g14291,g9839,g12155);
  NR2 NOR2_325(g11537,g8229,g3873);
  NR2 NOR2_326(g27343,g8005,g26616);
  NR2 NOR2_327(g28981,g9234,g27999);
  NR2 NOR2_328(g29077,g6555,g26994);
  NR2 NOR2_329(g12646,g9234,g9206);
  NR3 NOR3_27(g11283,g7953,g4991,g9064);
  NR2 NOR2_330(g10760,g1046,g7479);
  NR2 NOR2_331(g11303,g8497,g8500);
  NR2 NOR2_332(g31942,g8977,g30583);
  NR2 NOR2_333(g27368,g8119,g26657);
  NR2 NOR2_334(g21206,g6419,g17396);
  NR2 NOR2_335(g12850,g10430,g6845);
  NR2 NOR2_336(g13796,g9158,g12527);
  NR2 NOR2_337(g28521,g27649,g26604);
  NR2 NOR2_338(g31965,g30583,g4358);
  NR2 NOR2_339(g33131,g4659,g32057);
  NR4 NOR4_3(g12228,g10222,g10206,g10184,g10335);
  NR2 NOR2_340(g10649,g1183,g8407);
  NR3 NOR3_28(g12716,g7812,g6555,g6549);
  NR2 NOR2_341(g15123,g6975,g13605);
  NR2 NOR2_342(g10491,g6573,g9576);
  NR2 NOR2_343(g20027,g16242,g13779);
  NR2 NOR2_344(g21652,g17619,g17663);
  NR2 NOR2_345(g27379,g8492,g26636);
  NR2 NOR2_346(g11483,g8165,g3522);
  NR2 NOR2_347(g31469,g8822,g29725);
  NR2 NOR2_348(g11862,g7134,g7150);
  NR2 NOR2_349(g12050,g10038,g9649);
  NR2 NOR2_350(g24779,g3736,g23167);
  NR2 NOR2_351(g16237,g8088,g13574);
  NR3 NOR3_29(g29916,g8681,g28504,g11083);
  NR2 NOR2_352(g23135,g16476,g19981);
  NR2 NOR2_353(g15992,g10929,g13846);
  NR2 NOR2_354(g28462,g3512,g27617);
  NR2 NOR2_355(g13326,g10929,g10905);
  NR2 NOR2_356(g14767,g10130,g12204);
  NR2 NOR2_357(g14395,g12118,g9542);
  NR2 NOR2_358(g17420,g9456,g14408);
  NR2 NOR2_359(g10899,g4064,g8451);
  NR2 NOR2_360(g22540,g19720,g1373);
  NR2 NOR2_361(g11252,g8620,g3057);
  NR2 NOR2_362(g11621,g3512,g7985);
  NR2 NOR2_363(g15578,g7216,g14279);
  NR2 NOR2_364(g20998,g18065,g9450);
  NR2 NOR2_365(g33143,g32293,g31518);
  NR4 NOR4_4(g7661,g1211,g1216,g1221,g1205);
  NR2 NOR2_366(g29180,g9569,g26977);
  NR2 NOR2_367(g14247,g9934,g10869);
  NR2 NOR2_368(g13872,g8745,g11083);
  NR2 NOR2_369(g25501,g23918,g14645);
  NR2 NOR2_370(g20717,g5037,g17217);
  NR2 NOR2_371(g14272,g6411,g10598);
  NR2 NOR2_372(g12129,g9992,g7051);
  NR2 NOR2_373(g12002,g5297,g7004);
  NR3 NOR3_30(g11213,g4776,g7892,g9030);
  NR2 NOR2_374(g15142,g13680,g12889);
  NR2 NOR2_375(g33084,g31978,g7655);
  NR2 NOR2_376(g20149,g17091,g14185);
  NR2 NOR2_377(g26609,g146,g24732);
  NR2 NOR2_378(g15130,g13638,g6985);
  NR2 NOR2_379(g24148,g19268,g19338);
  NR2 NOR2_380(g15165,g12907,g13835);
  NR2 NOR2_381(g31373,g4975,g29725);
  NR2 NOR2_382(g11780,g4899,g8822);
  NR2 NOR2_383(g14360,g12078,g9484);
  NR2 NOR2_384(g9835,g2629,g2555);
  NR2 NOR2_385(g14447,g11938,g9698);
  NR2 NOR2_386(g12856,g10430,g6855);
  NR2 NOR2_387(g29187,g7704,g27999);
  NR3 NOR3_31(g11846,g7635,g7518,g7548);
  NR2 NOR2_388(g16209,g13478,g4749);
  NR2 NOR2_389(g14911,g10213,g12364);
  NR2 NOR2_390(g27499,g9095,g26636);
  NR3 NOR3_32(g28540,g8125,g27635,g7121);
  NR2 NOR2_391(g15372,g817,g14279);
  NR2 NOR2_392(g14754,g12821,g2988);
  NR2 NOR2_393(g27722,g7247,g25805);
  NR2 NOR2_394(g31117,g4991,g29556);
  NR2 NOR2_395(g27924,g9946,g25839);
  NR2 NOR2_396(g33117,g31261,g32205);
  NR2 NOR2_397(g22190,g2827,g18949);
  NR2 NOR2_398(g8720,g358,g365);
  NR2 NOR2_399(g15063,g6818,g13394);
  NR2 NOR2_400(g30934,g29836,g29850);
  NR2 NOR2_401(g19984,g17096,g8171);
  NR2 NOR2_402(g15137,g6992,g13680);
  NR2 NOR2_403(g12432,g1894,g8249);
  NR2 NOR2_404(g24959,g8858,g23324);
  NR2 NOR2_405(g17190,g723,g14279);
  NR2 NOR2_406(g14394,g12116,g9414);
  NR2 NOR2_407(g14367,g9547,g12289);
  NR2 NOR2_408(g16292,g7943,g13134);
  NR2 NOR2_409(g11357,g8558,g8561);
  NR3 NOR3_33(g29179,g9311,g28010,g7738);
  NR2 NOR2_410(g14420,g12153,g9490);
  NR2 NOR2_411(g12198,g9797,g9800);
  NR2 NOR2_412(g19853,g15746,g1052);
  NR3 NOR3_34(g27528,g8770,g26352,g11083);
  NR2 NOR2_413(g10318,g25,g22);
  NR2 NOR2_414(g14446,g12190,g9644);
  NR2 NOR2_415(g14227,g9863,g10838);
  NR2 NOR2_416(g20857,g17929,g9380);
  NR2 NOR2_417(g27960,g7134,g25791);
  NR2 NOR2_418(g14540,g12287,g9834);
  NR2 NOR2_419(g19401,g17193,g14296);
  NR2 NOR2_420(g17700,g14792,g12983);
  NR2 NOR2_421(g17625,g14541,g12123);
  NR2 NOR2_422(g15073,g12844,g13416);
  NR3 NOR3_35(g28481,g3506,g10323,g27617);
  NR2 NOR2_423(g10281,g5535,g5527);
  NR2 NOR2_424(g15122,g6959,g13605);
  NR2 NOR2_425(g26515,g24843,g24822);
  NR2 NOR2_426(g12708,g9518,g9462);
  NR2 NOR2_427(g25005,g6811,g23324);
  NR2 NOR2_428(g10699,g8526,g1514);
  NR2 NOR2_429(g15153,g13745,g12897);
  NR2 NOR2_430(g31116,g7892,g29540);
  NR3 NOR3_36(g11248,g7953,g4991,g4983);
  NR3 NOR3_37(g32780,g31327,I30330,I30331);
  NR2 NOR2_431(g15136,g13680,g12885);
  NR2 NOR2_432(g29908,g6918,g28471);
  NR2 NOR2_433(g27879,g9523,g25856);
  NR2 NOR2_434(g22450,g19345,g15724);
  NR3 NOR3_38(g12970,g10555,g10510,g10488);
  NR2 NOR2_435(g27878,g9559,g25839);
  NR2 NOR2_436(g27337,g8334,g26616);
  NR2 NOR2_437(g15164,g13835,g12906);
  NR2 NOR2_438(g11945,g7212,g7228);
  NR2 NOR2_439(g11999,g9654,g7423);
  NR2 NOR2_440(g10715,g8526,g8466);
  NR3 NOR3_39(g21389,g10143,g17748,g12259);
  NR2 NOR2_441(g20995,g5727,g17287);
  NR2 NOR2_442(g28520,g8229,g27635);
  NR2 NOR2_443(g25407,g23871,g14645);
  NR2 NOR2_444(g27010,g6052,g25839);
  NR2 NOR2_445(g11932,g843,g9166);
  NR2 NOR2_446(g33130,g32265,g31497);
  NR2 NOR2_447(g11448,g4191,g8790);
  NR2 NOR2_448(g14490,g9853,g12598);
  NR2 NOR2_449(g19907,g16210,g13676);
  NR2 NOR2_450(g21140,g6073,g17312);
  NR2 NOR2_451(g15091,g13177,g12863);
  NR2 NOR2_452(g33437,g31997,g10275);
  NR2 NOR2_453(g29007,g9269,g28010);
  NR2 NOR2_454(g10671,g1526,g8466);
  NR2 NOR2_455(g14181,g9083,g12259);
  NR2 NOR2_456(g23871,g2811,g21348);
  NR2 NOR2_457(g27353,g8097,g26616);
  NR2 NOR2_458(g16183,g9223,g13545);
  NR2 NOR2_459(g27823,g9792,g25805);
  NR4 NOR4_5(g11148,g8052,g9197,g9174,g9050);
  NR2 NOR2_460(g12680,g9631,g9576);
  NR2 NOR2_461(g19935,g17062,g8113);
  NR2 NOR2_462(g31372,g8796,g29697);
  NR2 NOR2_463(g25141,g22228,g10334);
  NR2 NOR2_464(g33175,g32099,g7828);
  NR2 NOR2_465(g24145,g19402,g19422);
  NR2 NOR2_466(g27966,g7153,g25805);
  NR3 NOR3_40(g13971,g8938,g4975,g11173);
  NR2 NOR2_467(g29035,g9321,g28020);
  NR2 NOR2_468(g14211,g9779,g10823);
  NR2 NOR2_469(g27364,g8426,g26616);
  NR2 NOR2_470(g33137,g4849,g32072);
  NR2 NOR2_471(g12017,g9969,g9586);
  NR2 NOR2_472(g12364,g10102,g10224);
  NR2 NOR2_473(g30613,g4507,g29365);
  NR2 NOR2_474(g29142,g5535,g28010);
  NR2 NOR2_475(g14497,g5990,g12705);
  NR2 NOR2_476(g30273,g5990,g29036);
  NR2 NOR2_477(g30106,g28739,g7268);
  NR2 NOR2_478(g12288,g2610,g8418);
  NR3 NOR3_41(g29193,g9529,g26994,g7812);
  NR2 NOR2_479(g19906,g16209,g13672);
  NR2 NOR2_480(g12571,g9511,g9451);
  NR2 NOR2_481(g12308,g9951,g9954);
  NR2 NOR2_482(g25004,g676,g23324);
  NR2 NOR2_483(g28496,g3179,g27602);
  NR2 NOR2_484(g29165,g5881,g28020);
  NR2 NOR2_485(g14339,g12289,g2735);
  NR2 NOR2_486(g16072,g10961,g13273);
  NR2 NOR2_487(g10338,g5062,g5022);
  NR2 NOR2_488(g15062,g6817,g13394);
  NR2 NOR2_489(g28986,g5517,g28010);
  NR2 NOR2_490(g29006,g5180,g27999);
  NR2 NOR2_491(g25947,g1199,g24591);
  NR2 NOR2_492(g15508,g10320,g14279);
  NR2 NOR2_493(g13959,g3698,g11309);
  NR2 NOR2_494(g27954,g10014,g25856);
  NR2 NOR2_495(g12752,g9576,g9529);
  NR2 NOR2_496(g11958,g9543,g7327);
  NR2 NOR2_497(g12374,g2185,g8205);
  NR2 NOR2_498(g13378,g11374,g11017);
  NR2 NOR2_499(g14411,g9460,g11160);
  NR2 NOR2_500(g13603,g8009,g10721);
  NR2 NOR2_501(g13944,g10262,g12259);
  NR2 NOR2_502(g14867,g10191,g12314);
  NR2 NOR2_503(g14450,g12195,g9598);
  NR2 NOR2_504(g29175,g6227,g26977);
  NR2 NOR2_505(g10819,g7479,g1041);
  NR2 NOR2_506(g13730,g3639,g11663);
  NR3 NOR3_42(g34359,g9162,g34174,g12259);
  NR2 NOR2_507(g14707,g10143,g12259);
  NR2 NOR2_508(g28457,g7980,g27602);
  NR3 NOR3_43(g32212,g8859,g31262,g11083);
  NR3 NOR3_44(g12558,g7738,g5517,g5511);
  NR2 NOR2_509(g13765,g8531,g11615);
  NR2 NOR2_510(g15051,g6801,g13350);
  NR2 NOR2_511(g15072,g13416,g12843);
  NR2 NOR2_512(g7192,g6444,g6404);
  NR2 NOR2_513(g29873,g6875,g28458);
  NR2 NOR2_514(g17180,g1559,g13574);
  NR3 NOR3_45(g22993,g1322,g16292,g19873);
  NR2 NOR2_515(g14094,g8770,g11083);
  NR2 NOR2_516(g15152,g13745,g12896);
  NR2 NOR2_517(g33109,g31997,g4584);
  NR2 NOR2_518(g12189,g1917,g8302);
  NR2 NOR2_519(g13129,g7553,g10762);
  NR2 NOR2_520(g10801,g1041,g7479);
  NR2 NOR2_521(g17694,g12435,g12955);
  NR2 NOR2_522(g33108,g32183,g31228);
  NR2 NOR2_523(g30134,g28768,g7280);
  NR3 NOR3_46(g11626,g7121,g3863,g3857);
  NR2 NOR2_524(g10695,g8462,g8407);
  NR2 NOR2_525(g27093,g26712,g26749);
  NR2 NOR2_526(g17619,g10179,g12955);
  NR2 NOR2_527(g12093,g9924,g7028);
  NR2 NOR2_528(g26649,g9037,g24732);
  NR2 NOR2_529(g27875,g9875,g25821);
  NR2 NOR2_530(g33174,g8714,g32072);
  NR3 NOR3_47(g11232,g4966,g7898,g9064);
  NR2 NOR2_531(g29034,g5527,g28010);
  NR2 NOR2_532(g19400,g17139,g14206);
  NR2 NOR2_533(g21127,g18065,g12099);
  NR2 NOR2_534(g11697,g8080,g3857);
  NR2 NOR2_535(g11995,g9645,g7410);
  NR2 NOR2_536(g16027,g10929,g13260);
  NR3 NOR3_48(g11261,g7928,g4801,g9030);
  NR2 NOR2_537(g14001,g739,g11083);
  NR2 NOR2_538(g30240,g7004,g28982);
  NR4 NOR4_6(g24631,g20516,g20436,g20219,g22957);
  NR2 NOR2_539(g12160,g9721,g9724);
  NR2 NOR2_540(g13512,g9077,g12527);
  NR2 NOR2_541(g28480,g8059,g27602);
  NR4 NOR4_7(g23956,g18957,g18918,g20136,g20114);
  NR2 NOR2_542(g8933,g4709,g4785);
  NR2 NOR2_543(g31483,g4899,g29725);
  NR2 NOR2_544(g13831,g11245,g7666);
  NR2 NOR2_545(g12201,g5417,g10047);
  NR2 NOR2_546(g29164,g9444,g28010);
  NR2 NOR2_547(g12467,g9472,g9407);
  NR2 NOR2_548(g30262,g5644,g29008);
  NR2 NOR2_549(g13989,g8697,g11309);
  NR2 NOR2_550(g13056,g7400,g10741);
  NR2 NOR2_551(g16090,g10961,g13315);
  NR2 NOR2_552(g26573,g24897,g24884);
  NR2 NOR2_553(g11924,g7187,g7209);
  NR2 NOR2_554(g29109,g9472,g26994);
  NR2 NOR2_555(g27352,g7975,g26616);
  NR2 NOR2_556(g26247,g7995,g24732);
  NR2 NOR2_557(g7781,g4064,g4057);
  NR2 NOR2_558(g12419,g9402,g9326);
  NR2 NOR2_559(g25770,g25417,g25377);
  NR2 NOR2_560(g29108,g6219,g26977);
  NR2 NOR2_561(g24976,g671,g23324);
  NR2 NOR2_562(g12418,g9999,g10001);
  NR2 NOR2_563(g12170,g10047,g5413);
  NR2 NOR2_564(g26098,g9073,g24732);
  NR2 NOR2_565(g23024,g7936,g19407);
  NR2 NOR2_566(g13342,g10961,g10935);
  NR2 NOR2_567(g13031,g7301,g10741);
  NR2 NOR2_568(g12853,g6848,g10430);
  NR3 NOR3_49(g33851,g8854,g33299,g12259);
  NR2 NOR2_569(g29174,g9511,g28020);
  NR3 NOR3_50(g21250,g9417,g9340,g17494);
  NR2 NOR2_570(g21658,g17694,g17727);
  NR2 NOR2_571(g22654,g7733,g19506);
  NR2 NOR2_572(g25521,g23955,g14645);
  NR3 NOR3_51(g11869,g7649,g7534,g7581);
  NR2 NOR2_573(g15647,g11924,g14248);
  NR2 NOR2_574(g28469,g3171,g27602);
  NR2 NOR2_575(g15090,g13144,g12862);
  NR3 NOR3_52(g28468,g3155,g10295,g27602);
  NR2 NOR2_576(g10341,g6227,g6219);
  NR2 NOR2_577(g25247,g23763,g14645);
  NR2 NOR2_578(g27704,g7239,g25791);
  NR2 NOR2_579(g11225,g3990,g6928);
  NR2 NOR2_580(g26162,g23052,g24751);
  NR3 NOR3_53(g16646,g13437,g11020,g11372);
  NR2 NOR2_581(g12466,g10057,g10059);
  NR2 NOR2_582(g25777,g25482,g25456);
  NR2 NOR2_583(g14335,g12045,g9283);
  NR2 NOR2_584(g12101,g6336,g7074);
  NR2 NOR2_585(g26628,g8990,g24732);
  NR2 NOR2_586(g29040,g6209,g26977);
  NR2 NOR2_587(g30162,g28880,g7462);
  NR2 NOR2_588(g8864,g3179,g3171);
  NR2 NOR2_589(g24383,g22409,g22360);
  NR2 NOR2_590(g27733,g9305,g25805);
  NR3 NOR3_54(g13970,g8883,g8796,g11155);
  NR4 NOR4_8(g11171,g8088,g9226,g9200,g9091);
  NR3 NOR3_55(g29183,g9392,g28020,g7766);
  NR3 NOR3_56(g24875,g8725,g23850,g11083);
  NR2 NOR2_591(g12166,g9856,g10124);
  NR3 NOR3_57(g14278,g562,g12259,g9217);
  NR2 NOR2_592(g13994,g4049,g11363);
  NR2 NOR2_593(g15149,g13745,g12894);
  NR2 NOR2_594(g25447,g23883,g14645);
  NR2 NOR2_595(g14306,g10060,g10887);
  NR3 NOR3_58(g29933,g8808,g28500,g12259);
  NR2 NOR2_596(g15148,g13716,g12893);
  NR2 NOR2_597(g15097,g12868,g13191);
  NR2 NOR2_598(g30147,g28768,g14567);
  NR2 NOR2_599(g13919,g3347,g11276);
  NR2 NOR2_600(g9755,g2070,g1996);
  NR2 NOR2_601(g13078,g7446,g10762);
  NR2 NOR2_602(g23695,g17420,g21140);
  NR2 NOR2_603(g19951,g16219,g13709);
  NR3 NOR3_59(g25776,g7166,g24380,g24369);
  NR2 NOR2_604(g25785,g25488,g25462);
  NR2 NOR2_605(g10884,g7650,g8451);
  NR2 NOR2_606(g27382,g8219,g26657);
  NR2 NOR2_607(g28953,g5170,g27999);
  NR2 NOR2_608(g24494,g23513,g23532);
  NR2 NOR2_609(g15133,g12883,g13638);
  NR3 NOR3_60(g32650,g31579,I30192,I30193);
  NR2 NOR2_610(g13125,g7863,g10762);
  NR2 NOR2_611(g10666,g8462,g1171);
  NR2 NOR2_612(g25950,g1070,g24591);
  NR2 NOR2_613(g7142,g6573,g6565);
  NR2 NOR2_614(g12154,g10155,g9835);
  NR2 NOR2_615(g29072,g9402,g26977);
  NR4 NOR4_9(g9602,g4688,g4681,g4674,g4646);
  NR2 NOR2_616(g14556,g6682,g12790);
  NR2 NOR2_617(g26645,g23602,g25160);
  NR2 NOR2_618(g13336,g11330,g11011);
  NR2 NOR2_619(g21256,g15483,g12179);
  NR3 NOR3_61(g22983,g979,g16268,g19853);
  NR2 NOR2_620(g9015,g3050,g3010);
  NR2 NOR2_621(g15050,g12834,g13350);
  NR2 NOR2_622(g12729,g1657,g8139);
  NR2 NOR2_623(g13631,g8068,g10733);
  NR2 NOR2_624(g10922,g7650,g4057);
  NR2 NOR2_625(g25446,g23686,g14645);
  NR2 NOR2_626(g22517,g19720,g1345);
  NR4 NOR4_10(g10179,g2098,g1964,g1830,g1696);
  NR4 NOR4_11(g9664,g4878,g4871,g4864,g4836);
  NR2 NOR2_627(g15096,g13191,g12867);
  NR2 NOR2_628(g30146,g28833,g7411);
  NR2 NOR2_629(g25540,g22409,g22360);
  NR2 NOR2_630(g14178,g8899,g11083);
  NR2 NOR2_631(g31482,g8883,g29697);
  NR2 NOR2_632(g30290,g6682,g29110);
  NR2 NOR2_633(g28568,g10323,g27617);
  NR2 NOR2_634(g25203,g6428,g23756);
  NR2 NOR2_635(g11309,g8587,g8728);
  NR3 NOR3_62(g11571,g10323,g3512,g3506);
  NR2 NOR2_636(g22523,g1345,g19720);
  NR2 NOR2_637(g14417,g12149,g9648);
  NR2 NOR2_638(g12622,g9569,g9518);
  NR2 NOR2_639(g26715,g23711,g25203);
  NR2 NOR2_640(g23763,g2795,g21276);
  NR2 NOR2_641(g14334,g12044,g9337);
  NR2 NOR2_642(g16232,g13516,g4950);
  NR2 NOR2_643(g11976,g9595,g7379);
  NR2 NOR2_644(g33090,g31997,g4593);
  NR3 NOR3_63(g31233,g8522,g29778,g24825);
  NR2 NOR2_645(g17727,g12486,g12983);
  NR2 NOR2_646(g11954,g9538,g7314);
  NR2 NOR2_647(g13954,g8663,g11276);
  NR2 NOR2_648(g28510,g3530,g27617);
  NR2 NOR2_649(g12333,g1624,g8139);
  NR2 NOR2_650(g26297,g8519,g24825);
  NR2 NOR2_651(g15129,g6984,g13638);
  NR2 NOR2_652(g12852,g6847,g10430);
  NR2 NOR2_653(g15057,g6810,g13350);
  NR2 NOR2_654(g11669,g3863,g8026);
  NR2 NOR2_655(g15128,g13638,g12880);
  NR2 NOR2_656(g14000,g8766,g12259);
  NR2 NOR2_657(g33449,g10311,g31950);
  NR2 NOR2_658(g33448,g7785,g31950);
  NR2 NOR2_659(g14568,g12000,g9915);
  NR2 NOR2_660(g17175,g1216,g13545);
  NR2 NOR2_661(g10123,g4294,g4297);
  NR2 NOR2_662(g21655,g17657,g17700);
  NR3 NOR3_64(g34354,g9003,g34162,g11083);
  NR3 NOR3_65(g12609,g7766,g5863,g5857);
  NR4 NOR4_12(g14751,g10622,g10617,g10609,g10603);
  NR2 NOR2_663(g14772,g6044,g12252);
  NR2 NOR2_664(g8182,g405,g392);
  NR2 NOR2_665(g28493,g3873,g27635);
  NR2 NOR2_666(g26546,g24858,g24846);
  NR2 NOR2_667(g19981,g3727,g16316);
  NR2 NOR2_668(g28340,g27439,g26339);
  NR2 NOR2_669(g14416,g12148,g9541);
  NR2 NOR2_670(g11610,g7980,g3155);
  NR2 NOR2_671(g25784,g25507,g25485);
  NR2 NOR2_672(g27973,g7187,g25839);
  NR2 NOR2_673(g33148,g4854,g32072);
  NR2 NOR2_674(g25956,g1413,g24609);
  NR2 NOR2_675(g11255,g8623,g6928);
  NR2 NOR2_676(g33097,g31950,g4628);
  NR2 NOR2_677(g14391,g12112,g9585);
  NR2 NOR2_678(g12798,g5535,g9381);
  NR3 NOR3_66(g10510,g7183,g4593,g4584);
  NR2 NOR2_679(g11270,g8431,g8434);
  NR2 NOR2_680(g16198,g9247,g13574);
  NR2 NOR2_681(g7352,g1526,g1514);
  NR2 NOR2_682(g26625,g23560,g25144);
  NR2 NOR2_683(g27732,g9364,g25791);
  NR3 NOR3_67(g13939,g4899,g8822,g11173);
  NR2 NOR2_684(g32017,g31504,g23475);
  NR2 NOR2_685(g26296,g8287,g24732);
  NR2 NOR2_686(g26338,g8458,g24825);
  NR2 NOR2_687(g15056,g6809,g13350);
  NR2 NOR2_688(g27400,g8553,g26657);
  NR2 NOR2_689(g10615,g1636,g7308);
  NR2 NOR2_690(g31133,g7953,g29556);
  NR2 NOR2_691(g33133,g32278,g31503);
  NR2 NOR2_692(g28475,g3863,g27635);
  NR2 NOR2_693(g21143,g15348,g9517);
  NR2 NOR2_694(g19388,g17181,g14256);
  NR2 NOR2_695(g15145,g12891,g13716);
  NR2 NOR2_696(g24439,g7400,g22312);
  NR2 NOR2_697(g9700,g2361,g2287);
  NR2 NOR2_698(g11201,g4125,g7765);
  NR2 NOR2_699(g33112,g31240,g32194);
  NR2 NOR2_700(g27771,g9809,g25839);
  NR2 NOR2_701(g19140,g7939,g15695);
  NR2 NOR2_702(g19997,g16231,g13739);
  NR2 NOR2_703(g15132,g12882,g13638);
  NR2 NOR2_704(g12235,g9234,g9206);
  NR2 NOR2_705(g33096,g31997,g4608);
  NR2 NOR2_706(g14362,g12080,g9338);
  NR2 NOR2_707(g22537,g19720,g1367);
  NR2 NOR2_708(g15161,g13809,g7073);
  NR2 NOR2_709(g14165,g8951,g11083);
  NR2 NOR2_710(g29104,g5188,g27999);
  NR2 NOR2_711(g12515,g9511,g5873);
  NR2 NOR2_712(g15087,g12860,g13144);
  NR2 NOR2_713(g32424,g8721,g31294);
  NR2 NOR2_714(g34496,g34370,g27648);
  NR2 NOR2_715(g14437,g9527,g11178);
  NR2 NOR2_716(g11194,g3288,g6875);
  NR2 NOR2_717(g15069,g6828,g13416);
  NR2 NOR2_718(g14347,g9309,g11123);
  NR3 NOR3_68(g14253,g10032,g12259,g9217);
  NR2 NOR2_719(g15068,g6826,g13416);
  NR2 NOR2_720(g17174,g9194,g14279);
  NR2 NOR2_721(g34067,g33859,g11772);
  NR2 NOR2_722(g11119,g9180,g9203);
  NR2 NOR2_723(g30150,g28846,g7424);
  NR2 NOR2_724(g33129,g8630,g32072);
  NR2 NOR2_725(g10821,g7503,g1384);
  NR4 NOR4_13(g12435,g9012,g8956,g8904,g8863);
  NR2 NOR2_726(g33128,g4653,g32057);
  NR2 NOR2_727(g14821,g6390,g12314);
  NR2 NOR2_728(g22522,g19699,g1024);
  NR2 NOR2_729(g11313,g8669,g3759);
  NR2 NOR2_730(g27345,g9360,g26636);
  NR2 NOR2_731(g12744,g9402,g6203);
  NR2 NOR2_732(g14516,g12227,g9704);
  NR2 NOR2_733(g11276,g8534,g8691);
  NR2 NOR2_734(g12849,g6840,g10430);
  NR2 NOR2_735(g17663,g10205,g12983);
  NR2 NOR2_736(g12848,g6839,g10430);
  NR2 NOR2_737(g27652,g3355,g26636);
  NR2 NOR2_738(g26256,g23873,g25479);
  NR2 NOR2_739(g22536,g1379,g19720);
  NR2 NOR2_740(g15086,g13144,g12859);
  NR2 NOR2_741(g12361,g6455,g10172);
  NR2 NOR2_742(g14726,g10090,g12166);
  NR2 NOR2_743(g30280,g7064,g29036);
  NR3 NOR3_69(g32455,g31566,I29985,I29986);
  NR2 NOR2_744(g15159,g13809,g12902);
  NR2 NOR2_745(g16288,g13794,g417);
  NR2 NOR2_746(g14320,g9257,g11111);
  NR2 NOR2_747(g15158,g13782,g12901);
  NR2 NOR2_748(g30157,g28833,g7369);
  NR2 NOR2_749(g14122,g8895,g12259);
  NR2 NOR2_750(g15144,g13716,g12890);
  NR2 NOR2_751(g31498,g9030,g29540);
  NR3 NOR3_70(g28492,g3857,g7121,g27635);
  NR3 NOR3_71(g8086,g168,g174,g182);
  NR2 NOR2_752(g11907,g7170,g7184);
  NR2 NOR2_753(g33432,g31997,g6978);
  NR2 NOR2_754(g26314,g24808,g24802);
  NR2 NOR2_755(g12371,g1760,g8195);
  NR2 NOR2_756(g23835,g2791,g21303);
  NR2 NOR2_757(g11238,g8584,g6905);
  NR2 NOR2_758(g17213,g11107,g13501);
  NR2 NOR2_759(g12234,g9776,g9778);
  NR2 NOR2_760(g23586,g17284,g20717);
  NR2 NOR2_761(g33145,g8677,g32072);
  NR2 NOR2_762(g14164,g9000,g12259);
  NR3 NOR3_72(g11185,g8038,g8183,g6804);
  NR2 NOR2_763(g13518,g3719,g11903);
  NR2 NOR2_764(g16488,g13697,g13656);
  NR2 NOR2_765(g16424,g8064,g13628);
  NR2 NOR2_766(g26268,g283,g24825);
  NR2 NOR2_767(g14575,g10050,g12749);
  NR2 NOR2_768(g11935,g9485,g7267);
  NR3 NOR3_73(g8131,g4776,g4801,g4793);
  NR2 NOR2_769(g27012,g6398,g25856);
  NR3 NOR3_74(g13883,g4709,g4785,g11155);
  NR2 NOR2_770(g33132,g4843,g32072);
  NR2 NOR2_771(g12163,g5073,g9989);
  NR2 NOR2_772(g28483,g8080,g27635);
  NR2 NOR2_773(g26993,g5360,g25805);
  NR2 NOR2_774(g33161,g32090,g7806);
  NR2 NOR2_775(g26667,g23642,g25175);
  NR2 NOR2_776(g30156,g28789,g14587);
  NR2 NOR2_777(g11729,g3179,g8059);
  NR2 NOR2_778(g13501,g3368,g11881);
  NR2 NOR2_779(g27829,g7345,g25856);
  NR2 NOR2_780(g14091,g8854,g12259);
  NR2 NOR2_781(g27828,g9892,g25856);
  NR3 NOR3_75(g22405,g18957,g20136,g20114);
  NR2 NOR2_782(g15669,g11945,g14272);
  NR2 NOR2_783(g12358,g10019,g10022);
  NR2 NOR2_784(g27344,g8390,g26636);
  NR2 NOR2_785(g12121,g10117,g9762);
  NR2 NOR2_786(g21193,g15348,g12135);
  NR2 NOR2_787(g22929,g19773,g12970);
  NR2 NOR2_788(g31068,g4801,g29540);
  NR2 NOR2_789(g11566,g3161,g7964);
  NR2 NOR2_790(g13622,g278,g11166);
  NR2 NOR2_791(g31970,g9024,g30583);
  NR2 NOR2_792(g12173,g10050,g7074);
  NR2 NOR2_793(g28509,g8107,g27602);
  NR2 NOR2_794(g16219,g13498,g4760);
  NR2 NOR2_795(g14522,g9924,g12656);
  NR2 NOR2_796(g11653,g7980,g7964);
  NR2 NOR2_797(g22357,g1024,g19699);
  NR3 NOR3_76(g29145,g6549,g7812,g26994);
  NR2 NOR2_798(g12029,g5644,g7028);
  NR2 NOR2_799(g10862,g7701,g7840);
  NR2 NOR2_800(g11415,g8080,g8026);
  NR2 NOR2_801(g29198,g7766,g28020);
  NR2 NOR2_802(g13852,g11320,g8347);
  NR2 NOR2_803(g30601,g16279,g29718);
  NR2 NOR2_804(g28452,g3161,g27602);
  NR2 NOR2_805(g27927,g9621,g25856);
  NR2 NOR2_806(g16201,g13462,g4704);
  NR2 NOR2_807(g15093,g13177,g6904);
  NR2 NOR2_808(g30143,g28761,g14566);
  NR2 NOR2_809(g23063,g16313,g19887);
  NR2 NOR2_810(g15065,g13394,g12840);
  NR2 NOR2_811(g30169,g28833,g14613);
  NR2 NOR2_812(g14397,g12120,g9416);
  NR2 NOR2_813(g12604,g5517,g9239);
  NR2 NOR2_814(g27770,g9386,g25821);
  NR2 NOR2_815(g19338,g16031,g1306);
  NR2 NOR2_816(g12755,g6555,g9407);
  NR2 NOR2_817(g33125,g8606,g32057);
  NR2 NOR2_818(g21209,g15483,g9575);
  NR2 NOR2_819(g14872,g6736,g12364);
  NR2 NOR2_820(g19968,g17062,g11223);
  NR2 NOR2_821(g23208,g20035,g16324);
  NR2 NOR2_822(g15160,g12903,g13809);
  NR2 NOR2_823(g13799,g8584,g11663);
  NR2 NOR2_824(g17482,g9523,g14434);
  NR2 NOR2_825(g33144,g4664,g32057);
  NR3 NOR3_77(g33823,g8774,g33306,g11083);
  NR2 NOR2_826(g20234,g17140,g14207);
  NR2 NOR2_827(g29069,g9381,g28010);
  NR2 NOR2_828(g11184,g513,g9040);
  NR2 NOR2_829(g7158,g5752,g5712);
  NR4 NOR4_14(g10205,g2657,g2523,g2389,g2255);
  NR2 NOR2_830(g24514,g23619,g23657);
  NR2 NOR2_831(g30922,g16662,g29810);
  NR2 NOR2_832(g29886,g3288,g28458);
  NR2 NOR2_833(g11692,g8021,g7985);
  NR2 NOR2_834(g16313,g8005,g13600);
  NR2 NOR2_835(g27926,g9467,g25856);
  NR2 NOR2_836(g13013,g7957,g10762);
  NR2 NOR2_837(g19070,g16957,g11720);
  NR2 NOR2_838(g22513,g1002,g19699);
  NR2 NOR2_839(g15155,g12899,g13782);
  NR2 NOR2_840(g11207,g3639,g6905);
  NR2 NOR2_841(g15170,g7118,g14279);
  NR2 NOR2_842(g22448,g1018,g19699);
  NR2 NOR2_843(g13539,g8594,g12735);
  NR2 NOR2_844(g13005,g7939,g10762);
  NR2 NOR2_845(g25321,g23835,g14645);
  NR2 NOR2_846(g14396,g12119,g9489);
  NR2 NOR2_847(g14731,g5698,g12204);
  NR2 NOR2_848(g15167,g13835,g12908);
  NR2 NOR2_849(g14413,g11914,g9638);
  NR2 NOR2_850(g28803,g27730,g22763);
  NR2 NOR2_851(g11771,g8921,g4185);
  NR2 NOR2_852(g25800,g25518,g25510);
  NR2 NOR2_853(g27766,g9716,g25791);
  NR2 NOR2_854(g23711,g9892,g21253);
  NR2 NOR2_855(g30117,g28739,g7252);
  NR2 NOR2_856(g29144,g9518,g26977);
  NR2 NOR2_857(g19402,g15979,g13133);
  NR2 NOR2_858(g23108,g16424,g19932);
  NR2 NOR2_859(g17148,g827,g14279);
  NR2 NOR2_860(g11414,g8591,g8593);
  NR2 NOR2_861(g16476,g8119,g13667);
  NR3 NOR3_78(g32585,g31542,I30123,I30124);
  NR2 NOR2_862(g15053,g12836,g13350);
  NR2 NOR2_863(g28482,g3522,g27617);
  NR2 NOR2_864(g30123,g28768,g7328);
  NR3 NOR3_79(g27629,g8891,g26382,g12259);
  NR2 NOR2_865(g28552,g10295,g27602);
  NR2 NOR2_866(g15101,g12871,g14591);
  NR2 NOR2_867(g12246,g9880,g9883);
  NR2 NOR2_868(g11584,g8229,g8172);
  NR2 NOR2_869(g30265,g7051,g29036);
  NR2 NOR2_870(g14640,g12371,g9824);
  NR2 NOR2_871(g15064,g6820,g13394);
  NR2 NOR2_872(g10803,g1384,g7503);
  NR2 NOR2_873(g12591,g504,g9040);
  NR2 NOR2_874(g12785,g9472,g6549);
  NR2 NOR2_875(g27355,g8443,g26657);
  NR2 NOR2_876(g13114,g7528,g10741);
  NR2 NOR2_877(g27825,g9316,g25821);
  NR2 NOR2_878(g11435,g8107,g3171);
  NR2 NOR2_879(g11107,g9095,g9177);
  NR2 NOR2_880(g15166,g13835,g7096);
  NR2 NOR2_881(g12858,g10365,g10430);
  NR2 NOR2_882(g11345,g8477,g8479);
  NR2 NOR2_883(g33093,g31997,g4601);
  NR2 NOR2_884(g31294,g11326,g29660);
  NR2 NOR2_885(g11940,g2712,g10084);
  NR2 NOR2_886(g27367,g8155,g26636);
  NR2 NOR2_887(g14027,g8734,g11363);
  NR2 NOR2_888(g11804,g8938,g4975);
  NR2 NOR2_889(g15570,g822,g14279);
  NR2 NOR2_890(g14248,g6065,g10578);
  NR2 NOR2_891(g16215,g1211,g13545);
  NR2 NOR2_892(g24990,g8898,g23324);
  NR2 NOR2_893(g14003,g9003,g11083);
  NR2 NOR2_894(g15074,g12845,g13416);
  NR2 NOR2_895(g12318,g10172,g6451);
  NR2 NOR2_896(g27059,g7577,g25895);
  NR3 NOR3_80(g15594,g10614,g13026,g7285);
  NR2 NOR2_897(g12059,g9853,g7004);
  NR2 NOR2_898(g12025,g9705,g7461);
  NR2 NOR2_899(g33160,g8672,g32057);
  NR2 NOR2_900(g12540,g2587,g8381);
  NR2 NOR2_901(g13500,g8480,g12641);
  NR2 NOR2_902(g15092,g12864,g13177);
  NR2 NOR2_903(g28149,g27598,g27612);
  NR2 NOR2_904(g15154,g13782,g12898);
  NR2 NOR2_905(g21062,g9547,g17297);
  NR2 NOR2_906(g14090,g8851,g12259);
  NR2 NOR2_907(g13004,g7933,g10741);
  NR2 NOR2_908(g33075,g31997,g7163);
  NR2 NOR2_909(g19268,g15979,g962);
  NR3 NOR3_81(g12377,g6856,g2748,g9708);
  NR2 NOR2_910(g12739,g9321,g9274);
  NR2 NOR2_911(g30130,g28761,g7275);
  NR3 NOR3_82(g24701,g979,g23024,g19778);
  NR2 NOR2_912(g12146,g1783,g8241);
  NR2 NOR2_913(g12645,g4467,g6961);
  NR2 NOR2_914(g13947,g8948,g11083);
  NR2 NOR2_915(g11273,g3061,g8620);
  NR2 NOR2_916(g14513,g12222,g9754);
  NR3 NOR3_83(g29705,g28399,g8284,g8404);
  NR2 NOR2_917(g14449,g12194,g9653);
  NR3 NOR3_84(g29189,g9462,g26977,g7791);
  NR2 NOR2_918(g33419,g31978,g7627);
  NR2 NOR2_919(g14448,g12192,g9699);
  NR2 NOR2_920(g11972,g9591,g7361);
  NR2 NOR2_921(g27366,g8016,g26636);
  NR2 NOR2_922(g7567,g979,g990);
  NR2 NOR2_923(g14212,g5373,g10537);
  NR2 NOR2_924(g12632,g9631,g6565);
  NR2 NOR2_925(g24766,g3385,g23132);
  NR2 NOR2_926(g23051,g7960,g19427);
  NR3 NOR3_85(g34703,g8899,g34545,g11083);
  NR3 NOR3_86(g11514,g10295,g3161,g3155);
  NR2 NOR2_927(g12226,g2476,g8373);
  NR2 NOR2_928(g31119,g7898,g29556);
  NR2 NOR2_929(g26873,g25374,g25331);
  NR2 NOR2_930(g11012,g7693,g7846);
  NR2 NOR2_931(g15139,g12886,g13680);
  NR2 NOR2_932(g26209,g23124,g24779);
  NR2 NOR2_933(g15138,g13680,g6993);
  NR2 NOR2_934(g11473,g8107,g8059);
  NR2 NOR2_935(g29915,g6941,g28484);
  NR2 NOR2_936(g27354,g8064,g26636);
  NR2 NOR2_937(g12297,g9269,g9239);
  NR2 NOR2_938(g13325,g7841,g10741);
  NR2 NOR2_939(g12980,g7909,g10741);
  NR2 NOR2_940(g12824,g5881,g9451);
  NR2 NOR2_941(g25952,g1542,g24609);
  NR2 NOR2_942(g13946,g8651,g11083);
  NR2 NOR2_943(g25175,g5736,g23692);
  NR2 NOR2_944(g14228,g5719,g10561);
  NR2 NOR2_945(g15585,g11862,g14194);
  NR2 NOR2_946(g26346,g8522,g24825);
  NR2 NOR2_947(g15608,g11885,g14212);
  NR2 NOR2_948(g15052,g12835,g13350);
  NR2 NOR2_949(g12211,g10099,g7097);
  NR2 NOR2_950(g31008,g30004,g30026);
  NR2 NOR2_951(g31476,g4709,g29697);
  NR2 NOR2_952(g29167,g9576,g26994);
  NR2 NOR2_953(g17198,g9282,g14279);
  NR2 NOR2_954(g27659,g3706,g26657);
  NR2 NOR2_955(g17393,g9386,g14379);
  NR2 NOR2_956(g12700,g9321,g5857);
  NR2 NOR2_957(g12659,g9451,g9392);
  NR2 NOR2_958(g12126,g9989,g5069);
  NR2 NOR2_959(g30136,g28799,g7380);
  NR2 NOR2_960(g19953,g16220,g13712);
  NR2 NOR2_961(g10793,g1389,g7503);
  NR2 NOR2_962(g14793,g2988,g12228);
  NR2 NOR2_963(g27338,g9291,g26616);
  NR2 NOR2_964(g12296,g9860,g9862);
  NR2 NOR2_965(g9762,g2495,g2421);
  NR2 NOR2_966(g23662,g17393,g20995);
  NR2 NOR2_967(g27969,g7170,g25821);
  NR2 NOR2_968(g14549,g9992,g12705);
  NR2 NOR2_969(g11755,g4709,g8796);
  NR2 NOR2_970(g29900,g3639,g28471);
  NR2 NOR2_971(g33092,g31978,g4332);
  NR2 NOR2_972(g11563,g8059,g8011);
  NR2 NOR2_973(g12855,g10430,g6854);
  NR2 NOR2_974(g31935,g30583,g4349);
  NR3 NOR3_87(g23204,g10685,g19462,g16488);
  NR2 NOR2_975(g14002,g8681,g11083);
  NR2 NOR2_976(g17657,g14751,g12955);
  NR3 NOR3_88(g11191,g4776,g4801,g9030);
  NR2 NOR2_977(g28498,g8172,g27635);
  NR2 NOR2_978(g15100,g13191,g12870);
  NR2 NOR2_979(g12581,g9569,g6219);
  NR2 NOR2_980(g33439,g31950,g4633);
  NR2 NOR2_981(g7175,g6098,g6058);
  NR2 NOR2_982(g33438,g31950,g4621);
  NR2 NOR2_983(g7139,g5406,g5366);
  NR2 NOR2_984(g22545,g1373,g19720);
  NR3 NOR3_89(g28031,g21209,I26522,I26523);
  NR2 NOR2_985(g12067,g5990,g7051);
  NR2 NOR2_986(g14512,g11955,g9753);
  NR2 NOR2_987(g27735,g7262,g25821);
  NR2 NOR2_988(g27877,g9397,g25839);
  NR3 NOR3_90(g28529,g8070,g27617,g10323);
  NR2 NOR2_989(g12150,g2208,g8259);
  NR2 NOR2_990(g33139,g8650,g32057);
  NR2 NOR2_991(g10831,g7690,g7827);
  NR2 NOR2_992(g13032,g7577,g10762);
  NR2 NOR2_993(g33138,g32287,g31514);
  NR2 NOR2_994(g14445,g12188,g9693);
  NR2 NOR2_995(g12695,g9269,g9239);
  NR3 NOR3_91(g29675,g28380,g8236,g8354);
  NR2 NOR2_996(g26183,g23079,g24766);
  NR2 NOR2_997(g30252,g7028,g29008);
  NR2 NOR2_998(g7304,g1183,g1171);
  NR2 NOR2_999(g14611,g12333,g9749);
  NR2 NOR2_1000(g7499,g333,g355);
  NR3 NOR3_92(g14988,g10816,g10812,g10805);
  NR2 NOR2_1001(g11360,g3763,g8669);
  NR2 NOR2_1002(g26872,g25411,g25371);
  NR2 NOR2_1003(g14271,g10002,g10874);
  NR2 NOR2_1004(g30183,g28880,g14644);
  NR2 NOR2_1005(g19430,g17150,g14220);
  NR2 NOR2_1006(g15141,g12888,g13680);
  NR2 NOR2_1007(g14145,g8945,g12259);
  NR2 NOR2_1008(g12256,g10136,g6105);
  NR2 NOR2_1009(g25948,g7752,g24609);
  NR2 NOR2_1010(g24497,g23533,g23553);
  NR2 NOR2_1011(g14529,g6336,g12749);
  NR2 NOR2_1012(g27102,g26750,g26779);
  NR2 NOR2_1013(g15135,g6990,g13638);
  NR2 NOR2_1014(g26574,g24887,g24861);
  NR2 NOR2_1015(g14393,g12115,g9488);
  NR2 NOR2_1016(g14365,g12084,g9339);
  NR3 NOR3_93(g32845,g30673,I30399,I30400);
  NR2 NOR2_1017(g17309,g9305,g14344);
  NR2 NOR2_1018(g15049,g13350,g6799);
  NR2 NOR2_1019(g11950,g9220,g9166);
  NR2 NOR2_1020(g10709,g7499,g351);
  NR3 NOR3_94(g27511,g22137,g26866,g20277);
  NR2 NOR2_1021(g12854,g6849,g10430);
  NR2 NOR2_1022(g28425,g27493,g26351);
  NR4 NOR4_15(g34912,g34883,g20277,g20242,g21370);
  NR3 NOR3_95(g25851,g4311,g24380,g24369);
  NR3 NOR3_96(g13996,g8938,g8822,g11173);
  NR3 NOR3_97(g28444,g8575,g27463,g24825);
  NR2 NOR2_1023(g15106,g12872,g10430);
  NR2 NOR2_1024(g17954,g832,g14279);
  NR2 NOR2_1025(g12550,g9300,g9259);
  NR2 NOR2_1026(g12314,g10053,g10207);
  NR2 NOR2_1027(g14602,g10099,g12790);
  NR2 NOR2_1028(g27721,g9672,g25805);
  NR2 NOR2_1029(g12085,g10082,g9700);
  NR2 NOR2_1030(g22488,g19699,g1002);
  NR2 NOR2_1031(g14337,g12049,g9284);
  NR3 NOR3_98(g11203,g4966,g4991,g9064);
  NR2 NOR2_1032(g13044,g7349,g10762);
  NR4 NOR4_16(g14792,g10653,g10623,g10618,g10611);
  NR3 NOR3_99(g28353,g9073,g27654,g24732);
  NR2 NOR2_1033(g29200,g7791,g26977);
  NR2 NOR2_1034(g9640,g1802,g1728);
  NR2 NOR2_1035(g19063,g7909,g15674);
  NR2 NOR2_1036(g33100,g32172,g31188);
  NR2 NOR2_1037(g13377,g7873,g10762);
  NR2 NOR2_1038(g14425,g5644,g12656);
  NR2 NOR2_1039(g27734,g9733,g25821);
  NR2 NOR2_1040(g15163,g13809,g12905);
  NR2 NOR2_1041(g30929,g29803,g29835);
  NR2 NOR2_1042(g19873,g15755,g1395);
  NR3 NOR3_100(g10918,g1532,g7751,g7778);
  NR2 NOR2_1043(g19422,g16031,g13141);
  NR2 NOR2_1044(g14444,g11936,g9692);
  NR3 NOR3_101(g12667,g7791,g6209,g6203);
  NR3 NOR3_102(g19209,g12971,g15614,g11320);
  NR3 NOR3_103(g13698,g528,g12527,g11185);
  NR2 NOR2_1045(g31515,g4983,g29556);
  NR2 NOR2_1046(g29184,g9631,g26994);
  NR2 NOR2_1047(g23626,g17309,g20854);
  NR2 NOR2_1048(g15724,g13858,g11374);
  NR2 NOR2_1049(g24018,I23162,I23163);
  NR2 NOR2_1050(g30282,g6336,g29073);
  NR2 NOR2_1051(g19453,g17199,g14316);
  NR2 NOR2_1052(g15121,g12874,g13605);
  NR2 NOR2_1053(g12443,g9374,g9300);
  NR2 NOR2_1054(g19436,g17176,g14233);
  NR2 NOR2_1055(g13661,g528,g11185);
  NR2 NOR2_1056(g11715,g8080,g8026);
  NR3 NOR3_104(g29005,g5164,g7704,g27999);
  NR2 NOR2_1057(g33107,g32180,g31223);
  NR2 NOR2_1058(g12601,g9381,g9311);
  NR2 NOR2_1059(g15134,g13638,g12884);
  NR2 NOR2_1060(g14364,g12083,g9415);
  NR2 NOR2_1061(g25769,g25453,g25414);
  NR2 NOR2_1062(g11385,g8021,g7985);

endmodule
