module s1494(VDD,CK,CLR,v0,v1,v13_D_10,v13_D_11,v13_D_12,v13_D_13,v13_D_14,
  v13_D_15,
  v13_D_16,v13_D_17,v13_D_18,v13_D_19,v13_D_20,v13_D_21,v13_D_22,v13_D_23,
  v13_D_24,v13_D_6,v13_D_7,v13_D_8,v13_D_9,v2,v3,v4,v5,v6);
input VDD,CK,CLR,v6,v5,v4,v3,v2,v1,v0;
output v13_D_24,v13_D_23,v13_D_22,v13_D_21,v13_D_20,v13_D_19,v13_D_18,v13_D_17,
  v13_D_16,v13_D_15,v13_D_14,v13_D_13,v13_D_12,v13_D_11,v13_D_10,v13_D_9,
  v13_D_8,v13_D_7,v13_D_6;

  wire v12,v13_D_5C,v11,v13_D_4C,v10,v13_D_3C,v9,v13_D_2C,v8,v13_D_1C,v7,
    v13_D_0C,v4E,C70DE,C70D,C104DE,C104D,C141DE,C141D,C191DE,C191D,C218DE,
    C218D,C180DE,C180D,C90DE,C90D,v3E,v1E,C30DE,C30D,C194DE,C194D,C117DE,C117D,
    C195DE,C195D,C208DE,C208D,C118DE,C118D,C138DE,C138D,C220DE,C220D,C166DE,
    C166D,C49DE,C49D,v5E,C81DE,C81D,C131DE,C131D,v0E,C144DE,C144D,C157DE,C157D,
    v11E,v6E,C129DE,C129D,v9E,v2E,v10E,v12E,C165DE,C165D,C83DE,C83D,C108DE,
    C108D,C124DE,C124D,v8E,v7E,II650,Av13_D_24B,II653,Av13_D_23B,II656,
    Av13_D_22B,II659,Av13_D_21B,II662,Av13_D_20B,II665,Av13_D_19B,II668,
    Av13_D_18B,II671,Av13_D_17B,II674,Av13_D_16B,II677,Av13_D_15B,II680,
    Av13_D_14B,II683,Av13_D_13B,II686,Av13_D_12B,II689,Av13_D_11B,II692,
    Av13_D_10B,II695,Av13_D_9B,II698,Av13_D_8B,II701,Av13_D_7B,II704,Av13_D_6B,
    II707,Av13_D_5B,v13_D_5,II710,Av13_D_4B,v13_D_4,II713,Av13_D_3B,v13_D_3,
    II716,Av13_D_2B,v13_D_2,II719,Av13_D_1B,v13_D_1,II722,Av13_D_0B,v13_D_0,
    IIII560,IIII559,IIII555,IIII554,IIII547,IIII546,IIII538,IIII537,IIII534,
    IIII533,IIII528,IIII524,IIII520,IIII518,IIII516,IIII514,II142,IIII513,
    IIII510,IIII508,IIII506,IIII505,IIII503,IIII501,IIII500,IIII498,IIII497,
    IIII495,IIII494,IIII492,IIII491,IIII489,IIII486,IIII485,IIII483,IIII482,
    IIII479,IIII478,IIII476,IIII475,IIII473,IIII471,IIII470,IIII468,IIII466,
    IIII464,IIII463,IIII461,IIII460,IIII457,IIII456,IIII453,IIII452,IIII450,
    IIII449,IIII447,IIII446,IIII444,IIII442,IIII441,IIII439,IIII438,IIII436,
    IIII435,IIII433,IIII432,IIII430,IIII429,IIII427,IIII425,IIII423,IIII420,
    IIII419,IIII417,IIII415,IIII414,IIII412,IIII409,IIII406,IIII405,II254,
    IIII403,IIII402,IIII399,IIII398,IIII396,IIII395,IIII393,IIII392,IIII390,
    IIII389,IIII387,IIII386,IIII384,IIII383,IIII381,IIII380,IIII378,IIII377,
    IIII375,C86D,IIII374,IIII372,IIII371,IIII369,IIII368,IIII366,IIII365,C56D,
    IIII363,C178D,IIII362,IIII360,C59D,IIII359,IIII357,IIII356,C50D,IIII354,
    IIII352,IIII350,IIII349,IIII347,IIII346,IIII344,IIII342,C159D,IIII341,
    IIII339,IIII338,IIII336,IIII335,IIII333,IIII332,II329,IIII329,IIII328,
    IIII326,IIII325,IIII323,C127D,IIII321,C33D,IIII320,IIII318,IIII317,IIII315,
    C155D,IIII314,IIII311,C71D,IIII310,IIII308,C111D,IIII306,IIII305,IIII303,
    C172D,IIII302,IIII300,C105D,IIII299,IIII297,C209D,IIII296,IIII294,C211D,
    II368,IIII293,IIII291,C142D,C213D,IIII288,C203D,IIII287,IIII285,C222D,
    IIII284,IIII282,C36D,IIII281,C29D,IIII280,C26D,IIII278,IIII276,C27D,
    IIII275,IIII273,C201D,IIII272,IIII270,C55D,IIII269,IIII267,C214D,IIII266,
    C200D,IIII263,C41D,IIII262,C42D,IIII260,C78D,IIII259,IIII257,C215D,IIII256,
    IIII254,C39D,IIII253,IIII251,IIII250,C77D,IIII248,C45D,IIII247,IIII245,
    C185D,IIII243,IIII242,C130D,IIII240,C125D,IIII239,IIII237,C221D,IIII236,
    C219D,IIII234,C167D,IIII233,C168D,IIII232,IIII230,C109D,IIII229,IIII227,
    C139D,IIII226,IIII224,C163D,IIII223,C160D,IIII222,C156D,IIII220,C51D,
    IIII219,IIII218,C44D,IIII216,C189D,IIII215,IIII213,C57D,IIII212,IIII210,
    C120D,IIII209,C119D,IIII208,C122D,IIII206,C150D,IIII205,IIII203,C34D,
    IIII202,IIII200,IIII199,C63D,IIII197,C158D,IIII196,C161D,IIII194,IIII192,
    IIII191,IIII189,IIII188,C175D,IIII186,IIII185,IIII183,C183D,IIII182,
    IIII180,C173D,IIII179,IIII177,C137D,IIII176,C145D,IIII175,IIII174,C143D,
    IIII173,C146D,IIII171,C193D,IIII170,IIII169,IIII167,IIII166,C205D,IIII164,
    C133D,IIII163,IIII161,IIII160,C65D,IIII158,C84D,IIII157,C82D,IIII156,C80D,
    IIII154,C40D,IIII153,C52D,IIII152,IIII151,IIII149,C112D,IIII148,IIII146,
    C223D,IIII145,C216D,IIII142,C169D,IIII141,C170D,IIII140,C210D,IIII137,C46D,
    IIII136,C47D,IIII134,C151D,IIII133,C152D,IIII131,IIII130,C60D,IIII129,C72D,
    IIII128,C69D,IIII127,C73D,IIII126,C58D,IIII124,C164D,IIII123,C162D,II548,
    C199D,IIII120,C123D,IIII119,C126D,IIII117,C35D,IIII116,C37D,IIII114,C97D,
    IIII113,C93D,IIII112,IIII111,C98D,IIII109,C179D,IIII108,C181D,IIII106,
    C114D,IIII105,C113D,IIII104,C107D,IIII103,C115D,IIII101,C128D,IIII100,
    C134D,IIII98,C87D,IIII97,C88D,IIII96,C85D,IIII95,C76D,IIII93,C147D,IIII92,
    C140D,IIII91,C148D,IIII89,C48D,IIII88,C43D,IIII87,C53D,IIII86,C54D,IIII84,
    C224D,IIII83,C225D,IIII82,C217D,IIII80,C192D,IIII79,IIII78,C196D,IIII76,
    C174D,IIII75,IIII73,C31D,IIII72,C38D,IIII71,C28D,IIII69,C202D,IIII68,C206D,
    IIII66,C100D,IIII65,IIII64,IIII63,C99D,IIII62,C95D,IIII60,C74D,IIII59,C67D,
    IIII58,C75D,C153D,IIII55,C187D,IIII54,C186D,IIII52,C135D,IIII51,C132D,
    IIII49,C176D,IIII48,C177D,IIII46,C110D,IIII45,C116D,IIII44,C106D,IIII43,
    IIII41,C96D,IIII40,C92D,IIII39,C103D,IIII38,C102D,IIII36,C89D,IIII35,C79D,
    IIII34,C91D,IIII32,C207D,II642,IIII31,IIII29,C190D,IIII28,C188D,IIII27,
    C184D,II491,II497,II542,II610;

  FD1 DFF_0(CK,v12,v13_D_5C);
  FD1 DFF_1(CK,v11,v13_D_4C);
  FD1 DFF_2(CK,v10,v13_D_3C);
  FD1 DFF_3(CK,v9,v13_D_2C);
  FD1 DFF_4(CK,v8,v13_D_1C);
  FD1 DFF_5(CK,v7,v13_D_0C);
  IV  NOT_0(v4E,v4);
  IV  NOT_1(C70DE,C70D);
  IV  NOT_2(C104DE,C104D);
  IV  NOT_3(C141DE,C141D);
  IV  NOT_4(C191DE,C191D);
  IV  NOT_5(C218DE,C218D);
  IV  NOT_6(C180DE,C180D);
  IV  NOT_7(C90DE,C90D);
  IV  NOT_8(v3E,v3);
  IV  NOT_9(v1E,v1);
  IV  NOT_10(C30DE,C30D);
  IV  NOT_11(C194DE,C194D);
  IV  NOT_12(C117DE,C117D);
  IV  NOT_13(C195DE,C195D);
  IV  NOT_14(C208DE,C208D);
  IV  NOT_15(C118DE,C118D);
  IV  NOT_16(C138DE,C138D);
  IV  NOT_17(C220DE,C220D);
  IV  NOT_18(C166DE,C166D);
  IV  NOT_19(C49DE,C49D);
  IV  NOT_20(v5E,v5);
  IV  NOT_21(C81DE,C81D);
  IV  NOT_22(C131DE,C131D);
  IV  NOT_23(v0E,v0);
  IV  NOT_24(C144DE,C144D);
  IV  NOT_25(C157DE,C157D);
  IV  NOT_26(v11E,v11);
  IV  NOT_27(v6E,v6);
  IV  NOT_28(C129DE,C129D);
  IV  NOT_29(v9E,v9);
  IV  NOT_30(v2E,v2);
  IV  NOT_31(v10E,v10);
  IV  NOT_32(v12E,v12);
  IV  NOT_33(C165DE,C165D);
  IV  NOT_34(C83DE,C83D);
  IV  NOT_35(C108DE,C108D);
  IV  NOT_36(C124DE,C124D);
  IV  NOT_37(v8E,v8);
  IV  NOT_38(v7E,v7);
  IV  NOT_39(II650,Av13_D_24B);
  IV  NOT_40(v13_D_24,II650);
  IV  NOT_41(II653,Av13_D_23B);
  IV  NOT_42(v13_D_23,II653);
  IV  NOT_43(II656,Av13_D_22B);
  IV  NOT_44(v13_D_22,II656);
  IV  NOT_45(II659,Av13_D_21B);
  IV  NOT_46(v13_D_21,II659);
  IV  NOT_47(II662,Av13_D_20B);
  IV  NOT_48(v13_D_20,II662);
  IV  NOT_49(II665,Av13_D_19B);
  IV  NOT_50(v13_D_19,II665);
  IV  NOT_51(II668,Av13_D_18B);
  IV  NOT_52(v13_D_18,II668);
  IV  NOT_53(II671,Av13_D_17B);
  IV  NOT_54(v13_D_17,II671);
  IV  NOT_55(II674,Av13_D_16B);
  IV  NOT_56(v13_D_16,II674);
  IV  NOT_57(II677,Av13_D_15B);
  IV  NOT_58(v13_D_15,II677);
  IV  NOT_59(II680,Av13_D_14B);
  IV  NOT_60(v13_D_14,II680);
  IV  NOT_61(II683,Av13_D_13B);
  IV  NOT_62(v13_D_13,II683);
  IV  NOT_63(II686,Av13_D_12B);
  IV  NOT_64(v13_D_12,II686);
  IV  NOT_65(II689,Av13_D_11B);
  IV  NOT_66(v13_D_11,II689);
  IV  NOT_67(II692,Av13_D_10B);
  IV  NOT_68(v13_D_10,II692);
  IV  NOT_69(II695,Av13_D_9B);
  IV  NOT_70(v13_D_9,II695);
  IV  NOT_71(II698,Av13_D_8B);
  IV  NOT_72(v13_D_8,II698);
  IV  NOT_73(II701,Av13_D_7B);
  IV  NOT_74(v13_D_7,II701);
  IV  NOT_75(II704,Av13_D_6B);
  IV  NOT_76(v13_D_6,II704);
  IV  NOT_77(II707,Av13_D_5B);
  IV  NOT_78(v13_D_5,II707);
  IV  NOT_79(II710,Av13_D_4B);
  IV  NOT_80(v13_D_4,II710);
  IV  NOT_81(II713,Av13_D_3B);
  IV  NOT_82(v13_D_3,II713);
  IV  NOT_83(II716,Av13_D_2B);
  IV  NOT_84(v13_D_2,II716);
  IV  NOT_85(II719,Av13_D_1B);
  IV  NOT_86(v13_D_1,II719);
  IV  NOT_87(II722,Av13_D_0B);
  IV  NOT_88(v13_D_0,II722);
  AN2 AND2_0(v13_D_5C,v13_D_5,CLR);
  AN2 AND2_1(v13_D_4C,v13_D_4,CLR);
  AN2 AND2_2(v13_D_3C,v13_D_3,CLR);
  AN2 AND2_3(v13_D_2C,v13_D_2,CLR);
  AN2 AND2_4(v13_D_1C,v13_D_1,CLR);
  AN2 AND2_5(v13_D_0C,v13_D_0,CLR);
  AN2 AND2_6(IIII560,v7E,v12E);
  AN2 AND2_7(IIII559,v8,v11);
  AN3 AND3_0(IIII555,v0,v8E,v11);
  AN3 AND3_1(IIII554,v2E,v8,v9E);
  AN2 AND2_8(IIII547,v10,v11E);
  AN2 AND2_9(IIII546,v0,v11);
  AN2 AND2_10(IIII538,v8,v12E);
  AN4 AND4_0(IIII537,v6E,v7E,v8E,v12);
  AN2 AND2_11(IIII534,v8E,v10E);
  AN2 AND2_12(IIII533,v9,v10);
  AN2 AND2_13(IIII528,v9E,v11);
  AN2 AND2_14(IIII524,v6,v11E);
  AN2 AND2_15(IIII520,v3E,v6E);
  AN2 AND2_16(IIII518,v9,v10E);
  AN2 AND2_17(IIII516,v1,v12);
  AN4 AND4_1(IIII514,v2,v7,v9E,C138DE);
  AN3 AND3_2(II142,v7E,v9,v11E);
  AN3 AND3_3(IIII513,v12E,C166DE,II142);
  AN2 AND2_18(IIII510,v9,v10);
  AN2 AND2_19(IIII508,v9E,v11E);
  AN4 AND4_2(IIII506,v7E,v9,v10E,v12E);
  AN4 AND4_3(IIII505,v7,v8,C138DE,C191DE);
  AN2 AND2_20(IIII503,v9E,C30DE);
  AN2 AND2_21(IIII501,v8E,v11E);
  AN3 AND3_4(IIII500,v8,v11,C83DE);
  AN2 AND2_22(IIII498,v8,C117DE);
  AN3 AND3_5(IIII497,v8E,v9E,C194DE);
  AN3 AND3_6(IIII495,v9,v11,C131DE);
  AN3 AND3_7(IIII494,v8E,v10,C108DE);
  AN2 AND2_23(IIII492,v10,v11E);
  AN2 AND2_24(IIII491,v10E,C138DE);
  AN2 AND2_25(IIII489,v8E,v11);
  AN4 AND4_4(IIII486,v6E,v8E,v12,C129DE);
  AN3 AND3_8(IIII485,v6,C141DE,C220DE);
  AN4 AND4_5(IIII483,v8E,v9E,v11E,C83DE);
  AN2 AND2_26(IIII482,v2,C220DE);
  AN2 AND2_27(IIII479,v0,v11);
  AN2 AND2_28(IIII478,v10E,C83DE);
  AN4 AND4_6(IIII476,v8E,v9,v11E,v12E);
  AN3 AND3_9(IIII475,v2E,v8,C138DE);
  AN2 AND2_29(IIII473,v0E,C30DE);
  AN3 AND3_10(IIII471,v1,v10E,v12);
  AN3 AND3_11(IIII470,v8,v12E,C83DE);
  AN2 AND2_30(IIII468,v9,C83DE);
  AN3 AND3_12(IIII466,v8E,v11E,v12E);
  AN3 AND3_13(IIII464,v8E,v10E,v11);
  AN2 AND2_31(IIII463,C165DE,C191DE);
  AN3 AND3_14(IIII461,v8E,v9,v12);
  AN3 AND3_15(IIII460,v2E,v12E,C165DE);
  AN3 AND3_16(IIII457,v6,C124DE,C90DE);
  AN2 AND2_32(IIII456,v9,C30DE);
  AN3 AND3_17(IIII453,v8E,v10E,v12);
  AN2 AND2_33(IIII452,v12E,C220DE);
  AN4 AND4_7(IIII450,v3,v8,C138DE,C104DE);
  AN2 AND2_34(IIII449,C108DE,C83DE);
  AN4 AND4_8(IIII447,v8E,v9,v10E,v12E);
  AN2 AND2_35(IIII446,v11E,C90DE);
  AN2 AND2_36(IIII444,v3E,v9E);
  AN3 AND3_18(IIII442,v7E,v8E,v9E);
  AN2 AND2_37(IIII441,v11,C220DE);
  AN3 AND3_19(IIII439,v6,v12,C124DE);
  AN3 AND3_20(IIII438,v0,v10,C144DE);
  AN3 AND3_21(IIII436,v8E,v9,C144DE);
  AN2 AND2_38(IIII435,v12,C165DE);
  AN2 AND2_39(IIII433,v10,C144DE);
  AN2 AND2_40(IIII432,v7,C90DE);
  AN3 AND3_22(IIII430,v1E,v9,v10E);
  AN2 AND2_41(IIII429,v9E,C30DE);
  AN3 AND3_23(IIII427,v8E,v9,v10);
  AN2 AND2_42(IIII425,v8E,v10E);
  AN2 AND2_43(IIII423,v3E,C157DE);
  AN3 AND3_24(IIII420,v2E,v7,C131DE);
  AN4 AND4_9(IIII419,v5E,v7E,v8E,C30DE);
  AN3 AND3_25(IIII417,v5E,v11E,v12E);
  AN3 AND3_26(IIII415,v8E,v11E,v12E);
  AN2 AND2_44(IIII414,v6,C138DE);
  AN3 AND3_27(IIII412,v3,v10E,v12E);
  AN2 AND2_45(IIII409,v9,v11E);
  AN3 AND3_28(IIII406,v8,v11,C117DE);
  AN3 AND3_29(IIII405,v8E,v9E,C194DE);
  AN4 AND4_10(II254,v1,v6,v7E,v8E);
  AN4 AND4_11(IIII403,v9,v12E,C124DE,II254);
  AN3 AND3_30(IIII402,v8,v9E,C30DE);
  AN2 AND2_46(IIII399,v8,C141D);
  AN2 AND2_47(IIII398,v12E,C118DE);
  AN2 AND2_48(IIII396,v10E,v12E);
  AN2 AND2_49(IIII395,C157D,v9E);
  AN2 AND2_50(IIII393,v10E,v12E);
  AN2 AND2_51(IIII392,C81D,v11E);
  AN2 AND2_52(IIII390,C220D,v10E);
  AN3 AND3_31(IIII389,v8,v9,v10);
  AN3 AND3_32(IIII387,v8E,v9E,C124DE);
  AN4 AND4_12(IIII386,v0,C104D,v8,C30DE);
  AN2 AND2_53(IIII384,v10E,C138DE);
  AN2 AND2_54(IIII383,C70D,C141DE);
  AN2 AND2_55(IIII381,C166D,v11E);
  AN2 AND2_56(IIII380,v2,v11);
  AN4 AND4_13(IIII378,C218D,v5E,v9,v12E);
  AN3 AND3_33(IIII377,v7,v10,C90DE);
  AN2 AND2_57(IIII375,C86D,v10E);
  AN2 AND2_58(IIII374,v9E,C30DE);
  AN2 AND2_59(IIII372,C129D,v12E);
  AN2 AND2_60(IIII371,v10E,C90DE);
  AN2 AND2_61(IIII369,v9,C124DE);
  AN2 AND2_62(IIII368,C30D,C90DE);
  AN4 AND4_14(IIII366,v8E,v9,v11E,v12E);
  AN3 AND3_34(IIII365,C56D,v8,v11);
  AN2 AND2_63(IIII363,v1E,C178D);
  AN2 AND2_64(IIII362,v8,C138DE);
  AN2 AND2_65(IIII360,v3E,C59D);
  AN2 AND2_66(IIII359,v12E,C165DE);
  AN2 AND2_67(IIII357,v10,v11E);
  AN2 AND2_68(IIII356,C50D,v10E);
  AN2 AND2_69(IIII354,C191D,v11);
  AN2 AND2_70(IIII352,v8,C124D);
  AN2 AND2_71(IIII350,v11,C117D);
  AN2 AND2_72(IIII349,C118D,v11E);
  AN2 AND2_73(IIII347,C90D,v10E);
  AN2 AND2_74(IIII346,v12,C191DE);
  AN2 AND2_75(IIII344,C83D,v12E);
  AN2 AND2_76(IIII342,C159D,v8E);
  AN2 AND2_77(IIII341,v11E,C118DE);
  AN2 AND2_78(IIII339,v8E,C144DE);
  AN2 AND2_79(IIII338,C108D,C165DE);
  AN2 AND2_80(IIII336,C124D,v12);
  AN2 AND2_81(IIII335,v12E,C218DE);
  AN2 AND2_82(IIII333,v11E,v12E);
  AN2 AND2_83(IIII332,C138D,v9E);
  AN3 AND3_35(II329,v3,v7E,v10);
  AN4 AND4_15(Av13_D_20B,C138DE,C220DE,C104D,II329);
  AN3 AND3_36(IIII329,v9,v12,C30D);
  AN3 AND3_37(IIII328,v3,v12E,C124DE);
  AN2 AND2_84(IIII326,C81DE,C129D);
  AN2 AND2_85(IIII325,v10,C90DE);
  AN2 AND2_86(IIII323,v10E,C127D);
  AN3 AND3_38(IIII321,C33D,v11E,v12E);
  AN2 AND2_87(IIII320,v11,C141D);
  AN2 AND2_88(IIII318,v11,C118D);
  AN2 AND2_89(IIII317,v10,v11E);
  AN3 AND3_39(IIII315,C155D,v12E,C129D);
  AN2 AND2_90(IIII314,v10,C90DE);
  AN2 AND2_91(IIII311,C71D,v9E);
  AN4 AND4_16(IIII310,v6E,v9,v12E,C124DE);
  AN2 AND2_92(IIII308,C111D,C144DE);
  AN2 AND2_93(IIII306,C129DE,C138D);
  AN2 AND2_94(IIII305,v9,C49DE);
  AN2 AND2_95(IIII303,C172D,v12E);
  AN2 AND2_96(IIII302,v11E,C157DE);
  AN2 AND2_97(IIII300,v0E,C105D);
  AN2 AND2_98(IIII299,v11E,C108DE);
  AN3 AND3_40(IIII297,C209D,C208D,v11);
  AN4 AND4_17(IIII296,v8E,v9E,C124DE,C83DE);
  AN4 AND4_18(IIII294,C211D,v3,v7E,v11E);
  AN3 AND3_41(II368,v7,v8,v9E);
  AN3 AND3_42(IIII293,C138DE,C118DE,II368);
  AN2 AND2_99(IIII291,C142D,v11);
  AN4 AND4_19(Av13_D_21B,C213D,v7E,v10E,v12E);
  AN2 AND2_100(IIII288,v7E,C203D);
  AN2 AND2_101(IIII287,v9,v11);
  AN2 AND2_102(IIII285,C222D,v10E);
  AN2 AND2_103(IIII284,v11E,C157DE);
  AN2 AND2_104(IIII282,C36D,v12);
  AN2 AND2_105(IIII281,v3E,C29D);
  AN2 AND2_106(IIII280,v1E,C26D);
  AN2 AND2_107(IIII278,v10E,C138DE);
  AN4 AND4_20(IIII276,C27D,v7E,v9,v12E);
  AN3 AND3_43(IIII275,v7,v8,C90DE);
  AN2 AND2_108(IIII273,C201D,v8);
  AN2 AND2_109(IIII272,v10E,C144DE);
  AN2 AND2_110(IIII270,v1E,C55D);
  AN3 AND3_44(IIII269,v11E,C108DE,C83DE);
  AN3 AND3_45(IIII267,C214D,v7E,v10E);
  AN3 AND3_46(IIII266,v7,C49DE,C220DE);
  AN3 AND3_47(Av13_D_16B,C200D,v8,v10);
  AN3 AND3_48(IIII263,v7E,v11,C41D);
  AN2 AND2_111(IIII262,C42D,v8);
  AN2 AND2_112(IIII260,v3E,C78D);
  AN3 AND3_49(IIII259,v12E,C129DE,C83DE);
  AN2 AND2_113(IIII257,C215D,v9E);
  AN3 AND3_50(IIII256,v9,v10,C138DE);
  AN2 AND2_114(IIII254,C39D,v8E);
  AN3 AND3_51(IIII253,v1E,v10E,C138DE);
  AN3 AND3_52(IIII251,v6E,v11E,v12E);
  AN3 AND3_53(IIII250,C77D,v3,C138DE);
  AN2 AND2_115(IIII248,C45D,v10E);
  AN2 AND2_116(IIII247,v10,C144DE);
  AN2 AND2_117(IIII245,C185D,v8E);
  AN3 AND3_54(IIII243,C131D,v9,C144DE);
  AN2 AND2_118(IIII242,C130D,C165DE);
  AN2 AND2_119(IIII240,C125D,v9E);
  AN3 AND3_55(IIII239,v9,v12,C124DE);
  AN3 AND3_56(IIII237,v7,v12E,C221D);
  AN3 AND3_57(IIII236,v2E,v8,C219D);
  AN2 AND2_120(IIII234,v8,C167D);
  AN2 AND2_121(IIII233,C168D,v8E);
  AN2 AND2_122(IIII232,C165D,C83DE);
  AN2 AND2_123(IIII230,C109D,v10E);
  AN3 AND3_58(IIII229,v9,v10,C144DE);
  AN3 AND3_59(IIII227,C139D,v8,v10);
  AN3 AND3_60(IIII226,v8E,v10E,C144DE);
  AN3 AND3_61(IIII224,C163D,v8E,v11);
  AN3 AND3_62(IIII223,v7E,C160D,v9E);
  AN2 AND2_124(IIII222,C156D,C83DE);
  AN2 AND2_125(IIII220,C51D,v12);
  AN2 AND2_126(IIII219,C49D,v9);
  AN3 AND3_63(IIII218,v12E,C44D,C83DE);
  AN2 AND2_127(IIII216,C189D,v9E);
  AN3 AND3_64(IIII215,v1,v9,C144DE);
  AN2 AND2_128(IIII213,C57D,v10E);
  AN2 AND2_129(IIII212,v9E,C49DE);
  AN2 AND2_130(IIII210,v9,C120D);
  AN2 AND2_131(IIII209,v8,C119D);
  AN2 AND2_132(IIII208,C122D,v11E);
  AN2 AND2_133(IIII206,v7,C150D);
  AN2 AND2_134(IIII205,v8E,C30DE);
  AN2 AND2_135(IIII203,C34D,v9);
  AN4 AND4_21(IIII202,v9E,C144DE,C83DE,C194DE);
  AN2 AND2_136(IIII200,v12E,C124D);
  AN2 AND2_137(IIII199,v9E,C63D);
  AN3 AND3_65(IIII197,C158D,v7,v11E);
  AN2 AND2_138(IIII196,C161D,v11);
  AN3 AND3_66(IIII194,v3,v12,C77D);
  AN3 AND3_67(IIII192,v8E,v9E,C44D);
  AN3 AND3_68(IIII191,v8,v11,C117DE);
  AN2 AND2_139(IIII189,v7,v12E);
  AN2 AND2_140(IIII188,C175D,v11);
  AN3 AND3_69(IIII186,v8,v11,C117DE);
  AN2 AND2_141(IIII185,v8E,C195DE);
  AN2 AND2_142(IIII183,C183D,v8);
  AN3 AND3_70(IIII182,v8E,v10E,C144DE);
  AN2 AND2_143(IIII180,C173D,v9E);
  AN3 AND3_71(IIII179,v9,v10,C144DE);
  AN2 AND2_144(IIII177,C137D,C127D);
  AN2 AND2_145(IIII176,v10E,C145D);
  AN2 AND2_146(IIII175,v9,C144D);
  AN2 AND2_147(IIII174,v8E,C143D);
  AN2 AND2_148(IIII173,C146D,v11E);
  AN2 AND2_149(IIII171,v8,C193D);
  AN2 AND2_150(IIII170,v10,v11E);
  AN2 AND2_151(IIII169,C195D,v8E);
  AN3 AND3_72(IIII167,v8,v11,C129D);
  AN2 AND2_152(IIII166,C205D,v10);
  AN2 AND2_153(IIII164,C133D,v8E);
  AN3 AND3_73(IIII163,v11E,v12E,C118DE);
  AN2 AND2_154(IIII161,C144DE,C191D);
  AN2 AND2_155(IIII160,v8,C65D);
  AN2 AND2_156(IIII158,C84D,v10E);
  AN2 AND2_157(IIII157,C82D,v9E);
  AN2 AND2_158(IIII156,C80D,v9);
  AN2 AND2_159(IIII154,v2,C40D);
  AN2 AND2_160(IIII153,C52D,v8E);
  AN3 AND3_74(IIII152,v8,v12E,C129DE);
  AN2 AND2_161(IIII151,v9,C138DE);
  AN2 AND2_162(IIII149,C112D,v10);
  AN3 AND3_75(IIII148,v9,v10E,C144DE);
  AN3 AND3_76(IIII146,C223D,v8E,v9E);
  AN3 AND3_77(IIII145,C49DE,C166DE,C220DE);
  AN3 AND3_78(Av13_D_23B,C216D,v7E,v8E);
  AN2 AND2_163(IIII142,v7E,C169D);
  AN2 AND2_164(IIII141,C170D,v8);
  AN3 AND3_79(IIII140,v8E,v10E,C144DE);
  AN3 AND3_80(Av13_D_18B,C210D,v7E,v12E);
  AN2 AND2_165(IIII137,v8,C46D);
  AN2 AND2_166(IIII136,C47D,C144DE);
  AN3 AND3_81(IIII134,v7E,v10,C151D);
  AN2 AND2_167(IIII133,C152D,v9);
  AN3 AND3_82(IIII131,v9,v11E,C157DE);
  AN2 AND2_168(IIII130,C60D,C83D);
  AN2 AND2_169(IIII129,v8E,C72D);
  AN2 AND2_170(IIII128,v8,C69D);
  AN2 AND2_171(IIII127,C73D,v10E);
  AN2 AND2_172(IIII126,v2,C58D);
  AN2 AND2_173(IIII124,C164D,v12E);
  AN2 AND2_174(IIII123,v8,C162D);
  AN3 AND3_83(II548,C199D,v4,v5E);
  AN3 AND3_84(Av13_D_15B,v7E,v12E,II548);
  AN2 AND2_175(IIII120,v7E,C123D);
  AN2 AND2_176(IIII119,C126D,v8);
  AN2 AND2_177(IIII117,v8E,C35D);
  AN2 AND2_178(IIII116,C37D,v9);
  AN2 AND2_179(IIII114,v9,C97D);
  AN3 AND3_85(IIII113,v2E,v12E,C93D);
  AN2 AND2_180(IIII112,v11E,v12);
  AN2 AND2_181(IIII111,C98D,v10E);
  AN4 AND4_22(IIII109,C179D,v2,v8,v11);
  AN2 AND2_182(IIII108,C181D,C83DE);
  AN2 AND2_183(IIII106,v8E,C114D);
  AN2 AND2_184(IIII105,v8,C113D);
  AN3 AND3_86(IIII104,v3,C107D,v12);
  AN2 AND2_185(IIII103,C115D,v10);
  AN3 AND3_87(IIII101,C127D,C128D,v12E);
  AN2 AND2_186(IIII100,C134D,v9E);
  AN3 AND3_88(IIII98,v8E,v12,C87D);
  AN2 AND2_187(IIII97,C88D,v11E);
  AN2 AND2_188(IIII96,v8,C85D);
  AN2 AND2_189(IIII95,C76D,C81DE);
  AN2 AND2_190(IIII93,v7E,C147D);
  AN2 AND2_191(IIII92,v7,C140D);
  AN2 AND2_192(IIII91,C148D,C131DE);
  AN2 AND2_193(IIII89,v7,C48D);
  AN2 AND2_194(IIII88,v2E,C43D);
  AN2 AND2_195(IIII87,C53D,v7E);
  AN2 AND2_196(IIII86,C54D,C165DE);
  AN2 AND2_197(IIII84,v7E,C224D);
  AN2 AND2_198(IIII83,C225D,v11);
  AN3 AND3_89(IIII82,v0E,C217D,C108DE);
  AN3 AND3_90(IIII80,v7,v12E,C192D);
  AN2 AND2_199(IIII79,v8,C170D);
  AN2 AND2_200(IIII78,v7E,C196D);
  AN2 AND2_201(IIII76,v7E,C174D);
  AN2 AND2_202(IIII75,C129DE,C144DE);
  AN3 AND3_91(IIII73,v7,C31D,v8);
  AN2 AND2_203(IIII72,C38D,v7E);
  AN2 AND2_204(IIII71,v2E,C28D);
  AN2 AND2_205(IIII69,v7,C202D);
  AN2 AND2_206(IIII68,C206D,v12E);
  AN3 AND3_92(IIII66,v8E,v12E,C100D);
  AN2 AND2_207(IIII65,v9,C185D);
  AN2 AND2_208(IIII64,v11E,C157DE);
  AN2 AND2_209(IIII63,v8,C99D);
  AN2 AND2_210(IIII62,v6E,C95D);
  AN2 AND2_211(IIII60,v7E,C74D);
  AN2 AND2_212(IIII59,v7,C67D);
  AN2 AND2_213(IIII58,C75D,C129DE);
  AN2 AND2_214(Av13_D_9B,C153D,v12E);
  AN2 AND2_215(IIII55,C187D,v12E);
  AN2 AND2_216(IIII54,C186D,v9E);
  AN2 AND2_217(IIII52,C135D,v7E);
  AN2 AND2_218(IIII51,C132D,v7);
  AN2 AND2_219(IIII49,v8,C176D);
  AN2 AND2_220(IIII48,C177D,v8E);
  AN2 AND2_221(IIII46,v7,C110D);
  AN2 AND2_222(IIII45,C116D,v7E);
  AN2 AND2_223(IIII44,v2E,C106D);
  AN3 AND3_93(IIII43,v8,v10,C108DE);
  AN3 AND3_94(IIII41,v7,v12E,C96D);
  AN2 AND2_224(IIII40,v2,C92D);
  AN2 AND2_225(IIII39,C103D,v10E);
  AN2 AND2_226(IIII38,C102D,v7E);
  AN2 AND2_227(IIII36,v7E,C89D);
  AN4 AND4_23(IIII35,C79D,v7,v9,v12E);
  AN2 AND2_228(IIII34,C91D,C165DE);
  AN2 AND2_229(IIII32,C207D,v2);
  AN3 AND3_95(II642,v7E,v8E,C124DE);
  AN3 AND3_96(IIII31,C108DE,C83DE,II642);
  AN2 AND2_230(IIII29,C190D,v10);
  AN2 AND2_231(IIII28,v7E,C188D);
  AN2 AND2_232(IIII27,C184D,v7);
  OR2 OR2_0(C138D,v11E,v12E);
  OR2 OR2_1(C218D,v7E,v10);
  OR2 OR2_2(C131D,v8E,v10);
  OR2 OR2_3(C220D,v8E,v9E);
  OR2 OR2_4(C155D,v2,v7);
  OR2 OR2_5(C83D,v4E,v5E);
  OR2 OR2_6(C117D,v9E,v2);
  OR2 OR2_7(C178D,IIII559,IIII560);
  OR2 OR2_8(C70D,v0,v11E);
  OR2 OR2_9(C157D,v10E,v12E);
  OR2 OR2_10(C151D,IIII554,IIII555);
  OR2 OR2_11(C127D,v5E,v4);
  OR2 OR2_12(C142D,v0,v12);
  OR2 OR2_13(C166D,v3E,v6E);
  OR2 OR2_14(C165D,v8E,v11);
  OR2 OR2_15(C30D,v10E,v11E);
  OR2 OR2_16(C159D,IIII546,IIII547);
  OR2 OR2_17(C194D,v0,v10E);
  OR2 OR2_18(C193D,v2,v11E);
  OR2 OR2_19(C81D,v2E,v12);
  OR2 OR2_20(C124D,v10,v11);
  OR2 OR2_21(C208D,v5,v4);
  OR2 OR2_22(C191D,v10E,v9);
  OR2 OR2_23(C59D,IIII537,IIII538);
  OR2 OR2_24(C108D,v9,v12);
  OR2 OR2_25(C47D,IIII533,IIII534);
  OR2 OR2_26(C33D,v6E,v10);
  OR2 OR2_27(C104D,v1,v6E);
  OR2 OR2_28(C144D,v11E,v12);
  OR2 OR2_29(C145D,IIII528,v12);
  OR2 OR2_30(C90D,v9,v12E);
  OR2 OR2_31(C141D,v10E,v12);
  OR2 OR2_32(C86D,v9,IIII524);
  OR2 OR2_33(C118D,v2E,v10E);
  OR2 OR2_34(C129D,v9,v10);
  OR2 OR2_35(C50D,IIII520,v11);
  OR2 OR2_36(C179D,v10,IIII518);
  OR2 OR2_37(C56D,v9,IIII516);
  OR2 OR2_38(C200D,IIII513,IIII514);
  OR2 OR2_39(C36D,C165DE,v10E);
  OR2 OR2_40(C163D,C129DE,IIII510);
  OR2 OR2_41(C203D,C70DE,IIII508);
  OR2 OR2_42(C92D,IIII505,IIII506);
  OR2 OR2_43(C201D,IIII503,v12E);
  OR2 OR2_44(C27D,IIII500,IIII501);
  OR2 OR2_45(C209D,IIII497,IIII498);
  OR2 OR2_46(C60D,IIII494,IIII495);
  OR2 OR2_47(C185D,IIII491,IIII492);
  OR2 OR2_48(C137D,C117DE,IIII489);
  OR2 OR2_49(C45D,C90DE,v11E);
  OR2 OR2_50(C211D,IIII485,IIII486);
  OR2 OR2_51(C213D,IIII482,IIII483);
  OR2 OR2_52(C79D,C131DE,v11);
  OR2 OR2_53(C172D,IIII478,IIII479);
  OR2 OR2_54(C55D,IIII475,IIII476);
  OR2 OR2_55(C44D,IIII473,C124DE);
  OR2 OR2_56(C41D,IIII470,IIII471);
  OR2 OR2_57(C93D,C191DE,IIII468);
  OR2 OR2_58(C29D,C138DE,IIII466);
  OR2 OR2_59(C96D,IIII463,IIII464);
  OR2 OR2_60(C214D,IIII460,IIII461);
  OR2 OR2_61(C168D,C159D,v9);
  OR2 OR2_62(C114D,IIII456,IIII457);
  OR2 OR2_63(C170D,C124DE,v9E);
  OR2 OR2_64(C78D,IIII452,IIII453);
  OR2 OR2_65(C105D,IIII449,IIII450);
  OR2 OR2_66(C95D,IIII446,IIII447);
  OR2 OR2_67(C98D,C144D,IIII444);
  OR2 OR2_68(C156D,IIII441,IIII442);
  OR2 OR2_69(C215D,IIII438,IIII439);
  OR2 OR2_70(C103D,IIII435,IIII436);
  OR2 OR2_71(C42D,IIII432,IIII433);
  OR2 OR2_72(C100D,IIII429,IIII430);
  OR2 OR2_73(C76D,C131DE,IIII427);
  OR2 OR2_74(C120D,C144D,IIII425);
  OR2 OR2_75(C39D,IIII423,v9);
  OR2 OR2_76(C49D,C141D,v11);
  OR2 OR2_77(C217D,IIII419,IIII420);
  OR2 OR2_78(C222D,C138DE,IIII417);
  OR2 OR2_79(C26D,IIII414,IIII415);
  OR2 OR2_80(C54D,C90DE,IIII412);
  OR2 OR2_81(C77D,C104D,v0E);
  OR2 OR2_82(C148D,C90DE,IIII409);
  OR2 OR2_83(C180D,C194DE,v11E);
  OR2 OR2_84(C128D,IIII405,IIII406);
  OR2 OR2_85(C106D,IIII402,IIII403);
  OR2 OR2_86(C111D,C83DE,v2);
  OR2 OR2_87(C146D,IIII398,IIII399);
  OR2 OR2_88(C158D,IIII395,IIII396);
  OR2 OR2_89(C82D,IIII392,IIII393);
  OR2 OR2_90(C221D,IIII389,IIII390);
  OR2 OR2_91(C107D,IIII386,IIII387);
  OR2 OR2_92(C71D,IIII383,IIII384);
  OR2 OR2_93(C167D,IIII380,IIII381);
  OR2 OR2_94(C219D,IIII377,IIII378);
  OR2 OR2_95(C87D,IIII374,IIII375);
  OR2 OR2_96(C130D,IIII371,IIII372);
  OR2 OR2_97(C31D,IIII368,IIII369);
  OR2 OR2_98(C57D,IIII365,IIII366);
  OR2 OR2_99(C189D,IIII362,IIII363);
  OR2 OR2_100(C75D,IIII359,IIII360);
  OR2 OR2_101(C51D,IIII356,IIII357);
  OR2 OR2_102(C192D,v8,IIII354);
  OR2 OR2_103(C150D,C30DE,IIII352);
  OR3 OR3_0(C119D,IIII349,v12,IIII350);
  OR2 OR2_104(C91D,IIII346,IIII347);
  OR2 OR2_105(C84D,C138DE,IIII344);
  OR2 OR2_106(C160D,IIII341,IIII342);
  OR2 OR2_107(C109D,IIII338,IIII339);
  OR2 OR2_108(C125D,IIII335,IIII336);
  OR2 OR2_109(C139D,IIII332,IIII333);
  OR2 OR2_110(C69D,IIII328,IIII329);
  OR2 OR2_111(C175D,IIII325,IIII326);
  OR2 OR2_112(C122D,v12,IIII323);
  OR2 OR2_113(C34D,IIII320,IIII321);
  OR3 OR3_1(C63D,v12E,IIII317,IIII318);
  OR2 OR2_114(C161D,IIII314,IIII315);
  OR2 OR2_115(C195D,C180DE,v9);
  OR2 OR2_116(C72D,IIII310,IIII311);
  OR2 OR2_117(C112D,IIII308,v9E);
  OR2 OR2_118(C183D,IIII305,IIII306);
  OR2 OR2_119(C173D,IIII302,IIII303);
  OR2 OR2_120(C115D,IIII299,IIII300);
  OR2 OR2_121(C210D,IIII296,IIII297);
  OR2 OR2_122(Av13_D_19B,IIII293,IIII294);
  OR3 OR3_2(C143D,C49DE,v9,IIII291);
  OR2 OR2_123(C205D,IIII287,IIII288);
  OR2 OR2_124(C223D,IIII284,IIII285);
  OR3 OR3_3(C37D,IIII280,IIII281,IIII282);
  OR2 OR2_125(C133D,C49DE,IIII278);
  OR2 OR2_126(C28D,IIII275,IIII276);
  OR2 OR2_127(C202D,IIII272,IIII273);
  OR2 OR2_128(C73D,IIII269,IIII270);
  OR2 OR2_129(Av13_D_22B,IIII266,IIII267);
  OR2 OR2_130(C43D,IIII262,IIII263);
  OR2 OR2_131(C88D,IIII259,IIII260);
  OR2 OR2_132(C216D,IIII256,IIII257);
  OR2 OR2_133(C40D,IIII253,IIII254);
  OR2 OR2_134(C80D,IIII250,IIII251);
  OR2 OR2_135(C46D,IIII247,IIII248);
  OR2 OR2_136(C186D,C49DE,IIII245);
  OR2 OR2_137(C132D,IIII242,IIII243);
  OR2 OR2_138(C126D,IIII239,IIII240);
  OR2 OR2_139(C225D,IIII236,IIII237);
  OR4 OR4_0(C169D,IIII232,IIII233,v12,IIII234);
  OR2 OR2_140(C110D,IIII229,IIII230);
  OR2 OR2_141(C140D,IIII226,IIII227);
  OR3 OR3_4(C164D,IIII222,IIII223,IIII224);
  OR3 OR3_5(C52D,IIII218,IIII219,IIII220);
  OR2 OR2_142(C190D,IIII215,IIII216);
  OR2 OR2_143(C58D,IIII212,IIII213);
  OR4 OR4_1(C123D,C157DE,IIII208,IIII209,IIII210);
  OR2 OR2_144(C152D,IIII205,IIII206);
  OR2 OR2_145(C35D,IIII202,IIII203);
  OR2 OR2_146(C65D,IIII199,IIII200);
  OR2 OR2_147(C162D,IIII196,IIII197);
  OR2 OR2_148(C97D,v11E,IIII194);
  OR2 OR2_149(C199D,IIII191,IIII192);
  OR2 OR2_150(C176D,IIII188,IIII189);
  OR2 OR2_151(C181D,IIII185,IIII186);
  OR2 OR2_152(C184D,IIII182,IIII183);
  OR2 OR2_153(C174D,IIII179,IIII180);
  OR3 OR3_6(II491,IIII173,IIII174,IIII175);
  OR3 OR3_7(C147D,IIII176,IIII177,II491);
  OR3 OR3_8(II497,C208DE,C83DE,IIII169);
  OR4 OR4_2(C196D,IIII170,v12,IIII171,II497);
  OR2 OR2_154(C206D,IIII166,IIII167);
  OR2 OR2_155(C134D,IIII163,IIII164);
  OR2 OR2_156(C67D,IIII160,IIII161);
  OR3 OR3_9(C85D,IIII156,IIII157,IIII158);
  OR4 OR4_3(C53D,IIII151,IIII152,IIII153,IIII154);
  OR2 OR2_157(C113D,IIII148,IIII149);
  OR2 OR2_158(C224D,IIII145,IIII146);
  OR3 OR3_10(Av13_D_11B,IIII140,IIII141,IIII142);
  OR2 OR2_159(C48D,IIII136,IIII137);
  OR2 OR2_160(C153D,IIII133,IIII134);
  OR3 OR3_11(II542,IIII126,IIII127,IIII128);
  OR4 OR4_4(C74D,IIII129,IIII130,IIII131,II542);
  OR2 OR2_161(Av13_D_10B,IIII123,IIII124);
  OR2 OR2_162(Av13_D_6B,IIII119,IIII120);
  OR2 OR2_163(C38D,IIII116,IIII117);
  OR4 OR4_5(C99D,IIII111,IIII112,IIII113,IIII114);
  OR2 OR2_164(C187D,IIII108,IIII109);
  OR4 OR4_6(C116D,IIII103,IIII104,IIII105,IIII106);
  OR2 OR2_165(C135D,IIII100,IIII101);
  OR4 OR4_7(C89D,IIII95,IIII96,IIII97,IIII98);
  OR3 OR3_12(Av13_D_8B,IIII91,IIII92,IIII93);
  OR4 OR4_8(Av13_D_1B,IIII86,IIII87,IIII88,IIII89);
  OR3 OR3_13(Av13_D_24B,IIII82,IIII83,IIII84);
  OR3 OR3_14(Av13_D_14B,IIII78,IIII79,IIII80);
  OR2 OR2_166(C177D,IIII75,IIII76);
  OR3 OR3_15(Av13_D_0B,IIII71,IIII72,IIII73);
  OR2 OR2_167(C207D,IIII68,IIII69);
  OR3 OR3_16(II610,IIII62,IIII63,IIII64);
  OR3 OR3_17(C102D,IIII65,IIII66,II610);
  OR3 OR3_18(Av13_D_2B,IIII58,IIII59,IIII60);
  OR2 OR2_168(C188D,IIII54,IIII55);
  OR2 OR2_169(Av13_D_7B,IIII51,IIII52);
  OR2 OR2_170(Av13_D_12B,IIII48,IIII49);
  OR4 OR4_9(Av13_D_5B,IIII43,IIII44,IIII45,IIII46);
  OR4 OR4_10(Av13_D_4B,IIII38,IIII39,IIII40,IIII41);
  OR3 OR3_19(Av13_D_3B,IIII34,IIII35,IIII36);
  OR2 OR2_171(Av13_D_17B,IIII31,IIII32);
  OR3 OR3_20(Av13_D_13B,IIII27,IIII28,IIII29);

endmodule
