module s1238(VDD,CK,G0,G1,G10,G11,G12,G13,G2,G3,G4,G45,G5,G530,G532,G535,
  G537,G539,
  G542,G546,G547,G548,G549,G550,G551,G552,G6,G7,G8,G9);
input VDD,CK,G0,G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13;
output G549,G550,G551,G552,G542,G546,G547,G548,G530,G532,G535,G537,G45,G539;

  wire G29,G502,G30,G503,G31,G504,G32,G505,G33,G506,G34,G507,G35,G508,G36,G509,
    G37,G510,G38,G511,G39,G512,G40,G513,G41,G514,G42,G515,G43,G516,G44,G517,
    G518,G46,G519,G50,G49,G55,G54,G59,G58,G64,G63,G67,G70,G72,G71,G75,G74,G78,
    G77,G87,G86,G90,G89,G98,G97,G99,G123,G122,G125,G132,G135,G134,G140,G160,
    G161,G167,G168,G170,G171,G180,G181,G192,G193,G199,G200,G203,G204,G207,G208,
    G212,G213,G214,G215,G221,G222,G223,G224,G231,G232,G234,G235,G272,G271,G275,
    G274,G282,G281,G475,G57,G476,G477,G276,G478,G279,G479,G194,G480,G179,G481,
    G129,G482,G241,G483,G182,G484,G485,G486,G68,G487,G534,G488,G172,G489,G273,
    G490,G190,G491,G492,G62,G493,G544,G494,G173,G495,G496,G188,G497,G205,G498,
    G195,G499,G280,G500,G501,G156,G520,G521,G522,G524,G525,G526,G527,G528,G529,
    G531,G533,G536,G538,G540,G541,G543,G545,G554,G553,G81,G288,G240,G283,G219,
    G289,G119,G290,G117,G157,G291,G138,G155,G303,G120,G304,G52,G158,G306,G307,
    G104,G308,G151,G311,G178,G312,G315,G250,G251,G317,G159,G245,G321,G322,G105,
    G196,G323,G144,G324,G183,G327,G328,G102,G329,G150,G330,G248,G249,G331,G257,
    G336,G337,G270,G338,G202,G339,G209,G340,G341,G118,G342,G73,G197,G343,G147,
    G344,G111,G189,G346,G82,G347,G348,G349,G108,G351,G169,G352,G164,G353,G92,
    G163,G354,G357,G265,G358,G83,G359,G360,G106,G361,G362,G363,G364,G109,G365,
    G137,G366,G367,G126,G371,G267,G372,G116,G373,G376,G377,G56,G378,G379,G211,
    G380,G93,G382,G100,G383,G131,G385,G386,G85,G387,G388,G114,G392,G393,G127,
    G396,G76,G397,G101,G398,G94,G399,G65,G400,G277,G401,G110,G402,G154,G403,
    G176,G404,G218,G405,G174,G406,G410,G411,G48,G412,G413,G201,G414,G415,G146,
    G142,G165,G416,G61,G417,G418,G60,G422,G80,G423,G128,G424,G177,G425,G426,
    G162,G427,G95,G428,G227,G429,G51,G225,G430,G431,G432,G145,G153,G433,G91,
    G434,G216,G435,G236,G436,G437,G66,G229,G438,G133,G439,G175,G440,G441,G442,
    G121,G443,G47,G444,G445,G53,G446,G79,G447,G448,G139,G449,G88,G451,G187,
    G452,G184,G453,G186,G457,G107,G458,G459,G198,G460,G115,G461,G462,G463,G148,
    G467,G468,G124,G469,G470,G149,G471,G191,G103,G112,G472,G136,G473,G143,G474,
    G242,G141,G152,G244,G261,G269,G166,G284,G285,G286,G287,G292,G293,G294,G295,
    G296,G297,G298,G299,G300,G301,G302,G305,G309,G310,G313,G314,G316,G318,G319,
    G320,G325,G326,G332,G238,G333,G334,G335,G345,G226,G350,G355,G356,G368,G369,
    G239,G370,G374,G375,G381,G384,G389,G390,G391,G220,G394,G395,G407,G408,G409,
    G419,G420,G421,G228,G450,G454,G455,G206,G456,G464,G465,G210,G466,G260,G237,
    G264,G69,G233,G256,G84,G262,G96,G266,G217,G113,G268,G130,G263,G258,G259,
    G252,G253,G185,G230,G243,G246,G523,G254,G255,G278,G247;

  FD1 DFF_0(CK,G29,G502);
  FD1 DFF_1(CK,G30,G503);
  FD1 DFF_2(CK,G31,G504);
  FD1 DFF_3(CK,G32,G505);
  FD1 DFF_4(CK,G33,G506);
  FD1 DFF_5(CK,G34,G507);
  FD1 DFF_6(CK,G35,G508);
  FD1 DFF_7(CK,G36,G509);
  FD1 DFF_8(CK,G37,G510);
  FD1 DFF_9(CK,G38,G511);
  FD1 DFF_10(CK,G39,G512);
  FD1 DFF_11(CK,G40,G513);
  FD1 DFF_12(CK,G41,G514);
  FD1 DFF_13(CK,G42,G515);
  FD1 DFF_14(CK,G43,G516);
  FD1 DFF_15(CK,G44,G517);
  FD1 DFF_16(CK,G45,G518);
  FD1 DFF_17(CK,G46,G519);
  IV  NOT_0(G50,G49);
  IV  NOT_1(G55,G54);
  IV  NOT_2(G59,G58);
  IV  NOT_3(G64,G63);
  IV  NOT_4(G67,G44);
  IV  NOT_5(G70,G43);
  IV  NOT_6(G72,G71);
  IV  NOT_7(G75,G74);
  IV  NOT_8(G78,G77);
  IV  NOT_9(G87,G86);
  IV  NOT_10(G90,G89);
  IV  NOT_11(G98,G97);
  IV  NOT_12(G99,G29);
  IV  NOT_13(G123,G122);
  IV  NOT_14(G125,G40);
  IV  NOT_15(G132,G42);
  IV  NOT_16(G135,G134);
  IV  NOT_17(G140,G33);
  IV  NOT_18(G160,G161);
  IV  NOT_19(G167,G168);
  IV  NOT_20(G170,G171);
  IV  NOT_21(G180,G181);
  IV  NOT_22(G192,G193);
  IV  NOT_23(G199,G200);
  IV  NOT_24(G203,G204);
  IV  NOT_25(G207,G208);
  IV  NOT_26(G212,G213);
  IV  NOT_27(G214,G215);
  IV  NOT_28(G221,G222);
  IV  NOT_29(G223,G224);
  IV  NOT_30(G231,G232);
  IV  NOT_31(G234,G235);
  IV  NOT_32(G272,G271);
  IV  NOT_33(G275,G274);
  IV  NOT_34(G282,G281);
  IV  NOT_35(G475,G57);
  IV  NOT_36(G476,G30);
  IV  NOT_37(G477,G276);
  IV  NOT_38(G478,G279);
  IV  NOT_39(G479,G194);
  IV  NOT_40(G480,G179);
  IV  NOT_41(G481,G129);
  IV  NOT_42(G482,G241);
  IV  NOT_43(G483,G182);
  IV  NOT_44(G484,G30);
  IV  NOT_45(G485,G276);
  IV  NOT_46(G486,G68);
  IV  NOT_47(G487,G534);
  IV  NOT_48(G488,G172);
  IV  NOT_49(G489,G273);
  IV  NOT_50(G490,G190);
  IV  NOT_51(G491,G194);
  IV  NOT_52(G492,G62);
  IV  NOT_53(G493,G544);
  IV  NOT_54(G494,G173);
  IV  NOT_55(G495,G273);
  IV  NOT_56(G496,G188);
  IV  NOT_57(G497,G205);
  IV  NOT_58(G498,G195);
  IV  NOT_59(G499,G280);
  IV  NOT_60(G500,G173);
  IV  NOT_61(G501,G156);
  IV  NOT_62(G520,G0);
  IV  NOT_63(G521,G1);
  IV  NOT_64(G522,G2);
  IV  NOT_65(G524,G3);
  IV  NOT_66(G525,G526);
  IV  NOT_67(G527,G4);
  IV  NOT_68(G528,G5);
  IV  NOT_69(G529,G6);
  IV  NOT_70(G531,G7);
  IV  NOT_71(G533,G8);
  IV  NOT_72(G536,G9);
  IV  NOT_73(G538,G10);
  IV  NOT_74(G540,G11);
  IV  NOT_75(G541,G12);
  IV  NOT_76(G543,G13);
  IV  NOT_77(G545,G544);
  IV  NOT_78(G546,G41);
  IV  NOT_79(G554,G553);
  AN2 AND2_0(G81,G288,G240);
  AN2 AND2_1(G283,G122,G219);
  AN3 AND3_0(G289,G2,G119,G156);
  AN3 AND3_1(G290,G117,G135,G157);
  AN2 AND2_2(G291,G138,G155);
  AN2 AND2_3(G303,G5,G120);
  AN2 AND2_4(G304,G52,G158);
  AN2 AND2_5(G306,G524,G78);
  AN2 AND2_6(G307,G6,G104);
  AN2 AND2_7(G308,G5,G151);
  AN3 AND3_2(G311,G0,G178,G179);
  AN2 AND2_8(G312,G180,G182);
  AN2 AND2_9(G315,G250,G251);
  AN2 AND2_10(G317,G159,G245);
  AN2 AND2_11(G321,G90,G50);
  AN3 AND3_3(G322,G522,G105,G196);
  AN2 AND2_12(G323,G2,G144);
  AN2 AND2_13(G324,G522,G183);
  AN3 AND3_4(G327,G4,G39,G157);
  AN3 AND3_5(G328,G5,G102,G155);
  AN2 AND2_14(G329,G150,G156);
  AN2 AND2_15(G330,G248,G249);
  AN2 AND2_16(G331,G213,G257);
  AN2 AND2_17(G336,G1,G188);
  AN2 AND2_18(G337,G270,G167);
  AN2 AND2_19(G338,G202,G203);
  AN3 AND3_6(G339,G533,G199,G209);
  AN2 AND2_20(G340,G8,G270);
  AN2 AND2_21(G341,G531,G118);
  AN2 AND2_22(G342,G73,G197);
  AN3 AND3_7(G343,G2,G528,G147);
  AN3 AND3_8(G344,G111,G189,G195);
  AN2 AND2_23(G346,G2,G82);
  AN2 AND2_24(G347,G135,G178);
  AN3 AND3_9(G348,G1,G97,G55);
  AN2 AND2_25(G349,G6,G108);
  AN4 AND4_0(G351,G524,G169,G221,G234);
  AN4 AND4_1(G352,G8,G135,G37,G164);
  AN3 AND3_10(G353,G11,G92,G163);
  AN2 AND2_26(G354,G0,G214);
  AN2 AND2_27(G357,G265,G232);
  AN2 AND2_28(G358,G7,G83);
  AN2 AND2_29(G359,G6,G31);
  AN2 AND2_30(G360,G8,G106);
  AN2 AND2_31(G361,G6,G202);
  AN2 AND2_32(G362,G129,G77);
  AN2 AND2_33(G363,G77,G205);
  AN2 AND2_34(G364,G2,G109);
  AN3 AND3_11(G365,G282,G137,G156);
  AN2 AND2_35(G366,G125,G155);
  AN2 AND2_36(G367,G126,G157);
  AN3 AND3_12(G371,G161,G168,G267);
  AN3 AND3_13(G372,G116,G275,G155);
  AN2 AND2_37(G373,G34,G160);
  AN2 AND2_38(G376,G533,G75);
  AN2 AND2_39(G377,G90,G56);
  AN2 AND2_40(G378,G89,G50);
  AN2 AND2_41(G379,G9,G211);
  AN2 AND2_42(G380,G6,G93);
  AN3 AND3_14(G382,G9,G100,G34);
  AN2 AND2_43(G383,G131,G155);
  AN3 AND3_15(G385,G529,G7,G49);
  AN2 AND2_44(G386,G536,G85);
  AN3 AND3_16(G387,G6,G274,G75);
  AN2 AND2_45(G388,G11,G114);
  AN2 AND2_46(G392,G132,G155);
  AN2 AND2_47(G393,G127,G34);
  AN3 AND3_17(G396,G76,G272,G155);
  AN3 AND3_18(G397,G101,G98,G157);
  AN3 AND3_19(G398,G94,G156,G158);
  AN3 AND3_20(G399,G520,G1,G65);
  AN2 AND2_48(G400,G0,G277);
  AN3 AND3_21(G401,G2,G110,G155);
  AN2 AND2_49(G402,G154,G183);
  AN2 AND2_50(G403,G11,G176);
  AN2 AND2_51(G404,G4,G218);
  AN3 AND3_22(G405,G3,G174,G189);
  AN2 AND2_52(G406,G87,G172);
  AN2 AND2_53(G410,G1,G205);
  AN2 AND2_54(G411,G48,G59);
  AN2 AND2_55(G412,G3,G207);
  AN3 AND3_23(G413,G8,G197,G201);
  AN2 AND2_56(G414,G199,G36);
  AN4 AND4_2(G415,G2,G146,G142,G165);
  AN3 AND3_24(G416,G61,G167,G169);
  AN3 AND3_25(G417,G13,G282,G70);
  AN3 AND3_26(G418,G524,G60,G172);
  AN3 AND3_27(G422,G0,G80,G155);
  AN2 AND2_57(G423,G541,G128);
  AN3 AND3_28(G424,G78,G174,G177);
  AN2 AND2_58(G425,G146,G176);
  AN3 AND3_29(G426,G37,G162,G38);
  AN3 AND3_30(G427,G541,G95,G165);
  AN2 AND2_59(G428,G212,G227);
  AN2 AND2_60(G429,G51,G225);
  AN2 AND2_61(G430,G177,G196);
  AN2 AND2_62(G431,G524,G67);
  AN2 AND2_63(G432,G145,G153);
  AN2 AND2_64(G433,G91,G154);
  AN3 AND3_31(G434,G165,G216,G231);
  AN2 AND2_65(G435,G135,G236);
  AN2 AND2_66(G436,G123,G77);
  AN2 AND2_67(G437,G66,G229);
  AN3 AND3_32(G438,G8,G146,G133);
  AN2 AND2_68(G439,G174,G175);
  AN2 AND2_69(G440,G38,G234);
  AN2 AND2_70(G441,G0,G236);
  AN2 AND2_71(G442,G541,G121);
  AN2 AND2_72(G443,G47,G162);
  AN3 AND3_33(G444,G64,G78,G211);
  AN2 AND2_73(G445,G53,G225);
  AN2 AND2_74(G446,G524,G79);
  AN2 AND2_75(G447,G11,G175);
  AN2 AND2_76(G448,G139,G153);
  AN2 AND2_77(G449,G88,G154);
  AN3 AND3_34(G451,G541,G554,G187);
  AN2 AND2_78(G452,G526,G184);
  AN2 AND2_79(G453,G545,G186);
  AN3 AND3_35(G457,G4,G107,G135);
  AN2 AND2_80(G458,G528,G209);
  AN2 AND2_81(G459,G77,G198);
  AN3 AND3_36(G460,G2,G81,G115);
  AN2 AND2_82(G461,G529,G531);
  AN2 AND2_83(G462,G192,G538);
  AN2 AND2_84(G463,G521,G148);
  AN2 AND2_85(G467,G522,G198);
  AN2 AND2_86(G468,G527,G124);
  AN2 AND2_87(G469,G163,G3);
  AN2 AND2_88(G470,G528,G149);
  AN3 AND3_37(G471,G191,G103,G112);
  AN3 AND3_38(G472,G136,G9,G190);
  AN2 AND2_89(G473,G11,G143);
  AN2 AND2_90(G474,G242,G77);
  AN2 AND2_91(G511,G163,G164);
  OR2 OR2_0(G47,G440,G441);
  OR2 OR2_1(G60,G413,G414);
  OR2 OR2_2(G61,G405,G406);
  OR2 OR2_3(G73,G339,G340);
  OR2 OR2_4(G79,G444,G445);
  OR2 OR2_5(G88,G446,G447);
  OR2 OR2_6(G91,G430,G431);
  OR2 OR2_7(G92,G351,G352);
  OR3 OR3_0(G93,G376,G377,G378);
  OR2 OR2_8(G95,G424,G425);
  OR2 OR2_9(G105,G321,G273);
  OR2 OR2_10(G106,G358,G359);
  OR2 OR2_11(G108,G346,G347);
  OR2 OR2_12(G110,G399,G400);
  OR2 OR2_13(G114,G385,G386);
  OR3 OR3_1(G115,G457,G458,G459);
  OR2 OR2_14(G118,G337,G338);
  OR2 OR2_15(G121,G438,G439);
  OR2 OR2_16(G126,G363,G364);
  OR4 OR4_0(G128,G415,G416,G417,G418);
  OR2 OR2_17(G131,G379,G380);
  OR2 OR2_18(G133,G434,G435);
  OR2 OR2_19(G137,G348,G349);
  OR2 OR2_20(G139,G442,G443);
  OR2 OR2_21(G141,G353,G354);
  OR2 OR2_22(G142,G403,G404);
  OR2 OR2_23(G145,G426,G427);
  OR2 OR2_24(G146,G336,G170);
  OR2 OR2_25(G147,G341,G342);
  OR2 OR2_26(G149,G467,G468);
  OR2 OR2_27(G150,G303,G304);
  OR3 OR3_2(G152,G306,G307,G308);
  OR2 OR2_28(G193,G6,G30);
  OR2 OR2_29(G224,G533,G31);
  OR2 OR2_30(G242,G469,G470);
  OR2 OR2_31(G244,G371,G159);
  OR2 OR2_32(G261,G283,G528);
  OR2 OR2_33(G269,G362,G529);
  OR2 OR2_34(G279,G317,G166);
  OR3 OR3_3(G284,G528,G272,G281);
  OR2 OR2_35(G285,G5,G479);
  OR2 OR2_36(G286,G9,G540);
  OR2 OR2_37(G287,G522,G81);
  OR2 OR2_38(G288,G1,G528);
  OR2 OR2_39(G292,G538,G75);
  OR2 OR2_40(G293,G7,G540);
  OR3 OR3_4(G294,G1,G117,G281);
  OR2 OR2_41(G295,G122,G491);
  OR2 OR2_42(G296,G89,G484);
  OR2 OR2_43(G297,G64,G274);
  OR2 OR2_44(G298,G5,G497);
  OR2 OR2_45(G299,G123,G77);
  OR2 OR2_46(G300,G87,G97);
  OR2 OR2_47(G301,G122,G486);
  OR2 OR2_48(G302,G4,G529);
  OR2 OR2_49(G305,G524,G55);
  OR2 OR2_50(G309,G272,G5);
  OR2 OR2_51(G310,G522,G135);
  OR2 OR2_52(G313,G521,G475);
  OR2 OR2_53(G314,G527,G57);
  OR2 OR2_54(G316,G531,G536);
  OR3 OR3_5(G318,G6,G8,G232);
  OR2 OR2_55(G319,G529,G489);
  OR2 OR2_56(G320,G76,G272);
  OR3 OR3_6(G325,G7,G536,G222);
  OR2 OR2_57(G326,G533,G232);
  OR2 OR2_58(G332,G529,G238);
  OR2 OR2_59(G333,G528,G6);
  OR2 OR2_60(G334,G3,G4);
  OR2 OR2_61(G335,G1,G78);
  OR2 OR2_62(G345,G529,G226);
  OR2 OR2_63(G350,G6,G536);
  OR2 OR2_64(G355,G11,G116);
  OR2 OR2_65(G356,G6,G476);
  OR2 OR2_66(G368,G533,G536);
  OR2 OR2_67(G369,G540,G239);
  OR2 OR2_68(G370,G538,G11);
  OR2 OR2_69(G374,G536,G538);
  OR2 OR2_70(G375,G10,G540);
  OR2 OR2_71(G381,G7,G71);
  OR2 OR2_72(G384,G529,G71);
  OR2 OR2_73(G389,G9,G274);
  OR2 OR2_74(G390,G89,G50);
  OR2 OR2_75(G391,G74,G220);
  OR2 OR2_76(G394,G5,G58);
  OR2 OR2_77(G395,G4,G134);
  OR2 OR2_78(G407,G6,G117);
  OR2 OR2_79(G408,G529,G77);
  OR2 OR2_80(G409,G528,G55);
  OR2 OR2_81(G419,G3,G5);
  OR2 OR2_82(G420,G522,G59);
  OR3 OR3_7(G421,G521,G2,G228);
  OR2 OR2_83(G450,G12,G171);
  OR3 OR3_8(G454,G481,G122,G77);
  OR2 OR2_84(G455,G78,G206);
  OR2 OR2_85(G456,G520,G78);
  OR2 OR2_86(G464,G72,G536);
  OR2 OR2_87(G465,G524,G210);
  OR2 OR2_88(G466,G538,G71);
  OR2 OR2_89(G530,G401,G402);
  OR2 OR2_90(G532,G422,G423);
  OR2 OR2_91(G535,G432,G433);
  OR2 OR2_92(G537,G448,G449);
  OR3 OR3_9(G539,G451,G452,G453);
  OR2 OR2_93(G544,G343,G344);
  OR2 OR2_94(G547,G382,G383);
  OR2 OR2_95(G548,G392,G393);
  OR4 OR4_1(G549,G396,G397,G398,G477);
  OR4 OR4_2(G550,G289,G290,G291,G485);
  OR3 OR3_10(G551,G327,G328,G329);
  OR3 OR3_11(G552,G365,G366,G367);
  OR3 OR3_12(G553,G322,G323,G324);
  ND3 NAND3_0(G48,G407,G408,G409);
  ND2 NAND2_0(G49,G9,G538);
  ND2 NAND2_1(G51,G260,G237);
  ND3 NAND3_1(G52,G298,G299,G219);
  ND2 NAND2_2(G53,G264,G237);
  ND2 NAND2_3(G54,G4,G6);
  ND2 NAND2_4(G56,G374,G375);
  ND2 NAND2_5(G57,G0,G2);
  ND2 NAND2_6(G58,G1,G3);
  ND2 NAND2_7(G62,G534,G32);
  ND2 NAND2_8(G63,G75,G8);
  ND2 NAND2_9(G65,G527,G228);
  ND2 NAND2_10(G66,G129,G101);
  ND2 NAND2_11(G68,G302,G528);
  ND3 NAND3_2(G69,G419,G420,G233);
  ND2 NAND2_12(G71,G8,G10);
  ND2 NAND2_13(G74,G9,G11);
  ND2 NAND2_14(G76,G0,G3);
  ND2 NAND2_15(G77,G4,G528);
  ND3 NAND3_3(G80,G421,G226,G256);
  ND2 NAND2_16(G82,G334,G335);
  ND2 NAND2_17(G83,G355,G356);
  ND2 NAND2_18(G84,G369,G370);
  ND2 NAND2_19(G85,G384,G239);
  ND2 NAND2_20(G86,G55,G3);
  ND2 NAND2_21(G89,G531,G8);
  ND3 NAND3_4(G94,G261,G181,G262);
  ND2 NAND2_22(G96,G313,G314);
  ND2 NAND2_23(G97,G2,G5);
  ND2 NAND2_24(G100,G381,G220);
  ND2 NAND2_25(G101,G3,G4);
  ND3 NAND3_5(G102,G320,G266,G210);
  ND3 NAND3_6(G103,G529,G7,G30);
  ND3 NAND3_7(G104,G122,G238,G240);
  ND2 NAND2_26(G107,G456,G1);
  ND2 NAND2_27(G109,G269,G219);
  ND2 NAND2_28(G111,G213,G217);
  ND2 NAND2_29(G112,G8,G31);
  ND2 NAND2_30(G113,G389,G390);
  ND2 NAND2_31(G116,G6,G9);
  ND2 NAND2_32(G117,G2,G4);
  ND2 NAND2_33(G119,G284,G285);
  ND2 NAND2_34(G120,G294,G295);
  ND2 NAND2_35(G122,G522,G3);
  ND2 NAND2_36(G124,G0,G206);
  ND2 NAND2_37(G127,G391,G268);
  ND2 NAND2_38(G129,G527,G5);
  ND2 NAND2_39(G130,G466,G9);
  ND2 NAND2_40(G134,G3,G5);
  ND2 NAND2_41(G136,G222,G224);
  ND2 NAND2_42(G138,G465,G263);
  ND3 NAND3_8(G143,G258,G193,G259);
  ND3 NAND3_9(G144,G215,G252,G253);
  ND3 NAND3_10(G148,G454,G455,G0);
  ND2 NAND2_43(G151,G305,G200);
  ND2 NAND2_44(G159,G6,G155);
  ND2 NAND2_45(G161,G316,G72);
  ND2 NAND2_46(G166,G7,G50);
  ND2 NAND2_47(G168,G75,G221);
  ND2 NAND2_48(G171,G553,G187);
  ND2 NAND2_49(G181,G2,G78);
  ND2 NAND2_50(G185,G525,G184);
  ND2 NAND2_51(G200,G527,G529);
  ND2 NAND2_52(G204,G521,G87);
  ND2 NAND2_53(G206,G287,G524);
  ND2 NAND2_54(G208,G68,G229);
  ND2 NAND2_55(G210,G520,G272);
  ND2 NAND2_56(G213,G64,G275);
  ND3 NAND3_11(G215,G135,G55,G212);
  ND2 NAND2_57(G217,G50,G230);
  ND2 NAND2_58(G219,G524,G55);
  ND2 NAND2_59(G220,G7,G71);
  ND2 NAND2_60(G222,G533,G10);
  ND2 NAND2_61(G226,G527,G59);
  ND2 NAND2_62(G228,G524,G5);
  ND2 NAND2_63(G232,G536,G164);
  ND2 NAND2_64(G233,G522,G135);
  ND2 NAND2_65(G235,G6,G536);
  ND3 NAND3_12(G237,G10,G75,G201);
  ND2 NAND2_66(G238,G2,G524);
  ND2 NAND2_67(G239,G7,G533);
  ND2 NAND2_68(G240,G4,G134);
  ND3 NAND3_13(G243,G368,G275,G34);
  ND2 NAND2_69(G245,G8,G34);
  ND2 NAND2_70(G246,G544,G186);
  ND2 NAND2_71(G248,G529,G36);
  ND3 NAND3_14(G249,G11,G273,G201);
  ND2 NAND2_72(G250,G13,G523);
  ND2 NAND2_73(G251,G543,G32);
  ND4 NAND4_0(G252,G3,G11,G35,G216);
  ND2 NAND2_74(G253,G87,G218);
  ND2 NAND2_75(G254,G1,G152);
  ND3 NAND3_15(G255,G309,G2,G529);
  ND2 NAND2_76(G256,G4,G69);
  ND2 NAND2_77(G257,G538,G230);
  ND3 NAND3_16(G258,G464,G103,G223);
  ND2 NAND2_78(G259,G130,G225);
  ND3 NAND3_17(G260,G528,G529,G191);
  ND2 NAND2_79(G262,G527,G278);
  ND2 NAND2_80(G263,G0,G99);
  ND2 NAND2_81(G264,G227,G241);
  ND2 NAND2_82(G265,G531,G50);
  ND2 NAND2_83(G266,G524,G96);
  ND2 NAND2_84(G267,G536,G84);
  ND2 NAND2_85(G268,G11,G113);
  ND2 NAND2_86(G270,G345,G204);
  ND2 NAND2_87(G271,G1,G4);
  ND2 NAND2_88(G273,G325,G326);
  ND2 NAND2_89(G274,G7,G10);
  ND3 NAND3_18(G276,G3,G543,G140);
  ND3 NAND3_19(G277,G394,G395,G81);
  ND3 NAND3_20(G278,G332,G333,G134);
  ND2 NAND2_90(G280,G46,G247);
  ND2 NAND2_91(G281,G523,G534);
  ND2 NAND2_92(G503,G286,G538);
  ND2 NAND2_93(G504,G292,G293);
  ND3 NAND3_21(G505,G300,G301,G181);
  ND2 NAND2_94(G508,G318,G319);
  ND2 NAND2_95(G510,G350,G235);
  ND2 NAND2_96(G512,G310,G233);
  ND3 NAND3_22(G518,G450,G185,G246);
  ND3 NAND3_23(G523,G254,G255,G208);
  ND3 NAND3_24(G526,G1,G2,G141);
  ND3 NAND3_25(G534,G296,G297,G166);
  ND3 NAND3_26(G542,G243,G244,G279);
  NR2 NOR2_0(G153,G522,G540);
  NR2 NOR2_1(G154,G12,G488);
  NR2 NOR2_2(G155,G13,G480);
  NR2 NOR2_3(G156,G12,G543);
  NR2 NOR2_4(G157,G13,G483);
  NR2 NOR2_5(G158,G521,G281);
  NR3 NOR3_0(G162,G533,G185,G498);
  NR2 NOR2_6(G163,G0,G4);
  NR2 NOR2_7(G164,G531,G10);
  NR2 NOR2_8(G165,G524,G529);
  NR2 NOR2_9(G169,G5,G7);
  NR2 NOR2_10(G172,G2,G171);
  NR2 NOR2_11(G173,G5,G495);
  NR2 NOR2_12(G174,G1,G496);
  NR2 NOR2_13(G175,G86,G500);
  NR2 NOR2_14(G176,G4,G494);
  NR2 NOR2_15(G177,G357,G533);
  NR2 NOR2_16(G178,G521,G4);
  NR2 NOR2_17(G179,G541,G280);
  NR2 NOR2_18(G182,G12,G62);
  NR2 NOR2_19(G183,G330,G3);
  NR3 NOR3_1(G184,G541,G13,G499);
  NR2 NOR2_20(G186,G282,G501);
  NR2 NOR2_21(G187,G13,G492);
  NR3 NOR3_2(G188,G543,G493,G282);
  NR2 NOR2_22(G189,G522,G54);
  NR2 NOR2_23(G190,G7,G11);
  NR2 NOR2_24(G191,G9,G482);
  NR2 NOR2_25(G194,G281,G271);
  NR2 NOR2_26(G195,G521,G134);
  NR3 NOR3_3(G196,G5,G540,G86);
  NR2 NOR2_27(G197,G540,G232);
  NR2 NOR2_28(G198,G520,G3);
  NR2 NOR2_29(G201,G528,G54);
  NR2 NOR2_30(G202,G10,G63);
  NR2 NOR2_31(G205,G529,G122);
  NR2 NOR2_32(G209,G1,G524);
  NR2 NOR2_33(G211,G6,G274);
  NR2 NOR2_34(G216,G4,G5);
  NR2 NOR2_35(G218,G528,G217);
  NR2 NOR2_36(G225,G7,G8);
  NR2 NOR2_37(G227,G5,G200);
  NR2 NOR2_38(G229,G1,G522);
  NR2 NOR2_39(G230,G8,G490);
  NR3 NOR3_4(G236,G536,G274,G54);
  NR2 NOR2_40(G241,G10,G11);
  NR4 NOR4_0(G247,G471,G472,G473,G474);
  NR2 NOR2_41(G502,G436,G437);
  NR2 NOR2_42(G506,G311,G312);
  NR3 NOR3_5(G507,G315,G12,G487);
  NR2 NOR2_43(G509,G331,G5);
  NR2 NOR2_44(G513,G360,G361);
  NR3 NOR3_6(G514,G372,G373,G478);
  NR2 NOR2_45(G515,G387,G388);
  NR3 NOR3_7(G516,G410,G411,G412);
  NR2 NOR2_46(G517,G428,G429);
  NR4 NOR4_1(G519,G460,G461,G462,G463);

endmodule
