module s15850(VDD,CK,g100,g101,g102,g103,g10377,g10379,g104,g10455,g10457,
  g10459,
  g10461,g10463,g10465,g10628,g10801,g109,g11163,g11206,g11489,g1170,g1173,
  g1176,g1179,g1182,g1185,g1188,g1191,g1194,g1197,g1200,g1203,g1696,g1700,
  g1712,g18,g1957,g1960,g1961,g23,g2355,g2601,g2602,g2603,g2604,g2605,g2606,
  g2607,g2608,g2609,g2610,g2611,g2612,g2648,g27,g28,g29,g2986,g30,g3007,g3069,
  g31,g3327,g41,g4171,g4172,g4173,g4174,g4175,g4176,g4177,g4178,g4179,g4180,
  g4181,g4191,g4192,g4193,g4194,g4195,g4196,g4197,g4198,g4199,g42,g4200,g4201,
  g4202,g4203,g4204,g4205,g4206,g4207,g4208,g4209,g4210,g4211,g4212,g4213,
  g4214,g4215,g4216,g43,g44,g45,g46,g47,g48,g4887,g4888,g5101,g5105,g5658,
  g5659,g5816,g6253,g6254,g6255,g6256,g6257,g6258,g6259,g6260,g6261,g6262,
  g6263,g6264,g6265,g6266,g6267,g6268,g6269,g6270,g6271,g6272,g6273,g6274,
  g6275,g6276,g6277,g6278,g6279,g6280,g6281,g6282,g6283,g6284,g6285,g6842,
  g6920,g6926,g6932,g6942,g6949,g6955,g741,g742,g743,g744,g750,g7744,g8061,
  g8062,g82,g8271,g83,g8313,g8316,g8318,g8323,g8328,g8331,g8335,g8340,g8347,
  g8349,g8352,g84,g85,g8561,g8562,g8563,g8564,g8565,g8566,g86,g87,g872,g873,
  g877,g88,g881,g886,g889,g89,g892,g895,g8976,g8977,g8978,g8979,g898,g8980,
  g8981,g8982,g8983,g8984,g8985,g8986,g90,g901,g904,g907,g91,g910,g913,g916,
  g919,g92,g922,g925,g93,g94,g9451,g95,g96,g99,g9961);
input VDD,CK,g18,g27,g109,g741,g742,g743,g744,g872,g873,g877,g881,g1712,
  g1960,g1961,
  g1696,g750,g85,g42,g1700,g102,g104,g101,g29,g28,g103,g83,g23,g87,g922,g892,
  g84,g919,g1182,g925,g48,g895,g889,g1185,g41,g43,g99,g1173,g1203,g1188,g1197,
  g46,g31,g45,g92,g89,g898,g91,g93,g913,g82,g88,g1194,g47,g96,g910,g95,g904,
  g1176,g901,g44,g916,g100,g886,g30,g86,g1170,g1200,g1191,g907,g90,g94,g1179;
output g2355,g2601,g2602,g2603,g2604,g2605,g2606,g2607,g2608,g2609,g2610,g2611,
  g2612,g2648,g2986,g3007,g3069,g4172,g4173,g4174,g4175,g4176,g4177,g4178,
  g4179,g4180,g4181,g4887,g4888,g5101,g5105,g5658,g5659,g5816,g6920,g6926,
  g6932,g6942,g6949,g6955,g7744,g8061,g8062,g8271,g8313,g8316,g8318,g8323,
  g8328,g8331,g8335,g8340,g8347,g8349,g8352,g8561,g8562,g8563,g8564,g8565,
  g8566,g8976,g8977,g8978,g8979,g8980,g8981,g8982,g8983,g8984,g8985,g8986,
  g9451,g9961,g10377,g10379,g10455,g10457,g10459,g10461,g10463,g10465,g10628,
  g10801,g11163,g11206,g11489,g6842,g4171,g6267,g6257,g1957,g6282,g6284,g6281,
  g6253,g6285,g6283,g6265,g3327,g6269,g4204,g4193,g6266,g4203,g4212,g4196,
  g6263,g4194,g4192,g4213,g6256,g6258,g6279,g4209,g4208,g4214,g4206,g6261,
  g6255,g6260,g6274,g6271,g4195,g6273,g6275,g4201,g6264,g6270,g4216,g6262,
  g6278,g4200,g6277,g4198,g4210,g4197,g6259,g4202,g6280,g4191,g6254,g6268,
  g4205,g4207,g4215,g4199,g6272,g6276,g4211;

  wire g1289,g5660,g1882,g9349,g312,g5644,g452,g11257,g123,g8272,g207,g7315,
    g713,g9345,g1153,g6304,g1209,g10873,g1744,g5663,g1558,g7349,g695,g9343,
    g461,g11467,g940,g8572,g976,g11471,g709,g8432,g1092,g6810,g1574,g7354,
    g1864,g7816,g369,g11439,g1580,g7356,g1736,g6846,g39,g10774,g1651,g11182,
    g1424,g7330,g1737,g1672,g11037,g1077,g6805,g1231,g8279,g4,g8079,g774,g7785,
    g1104,g6815,g1304,g7290,g243,g7325,g1499,g8447,g1044,g7789,g1444,g8987,
    g757,g11179,g786,g8436,g1543,g7344,g552,g11045,g315,g5645,g1534,g7341,g622,
    g9338,g1927,g9354,g1660,g11033,g278,g7765,g1436,g8989,g718,g8433,g76,g7775,
    g554,g11047,g496,g11333,g981,g11472,g878,g4896,g590,g5653,g829,g4182,g1095,
    g6811,g704,g9344,g1265,g7302,g1786,g7814,g682,g8429,g1296,g7292,g587,g6295,
    g52,g7777,g646,g8065,g327,g5649,g1389,g6836,g1371,g7311,g1956,g1955,g1675,
    g11038,g354,g11508,g113,g7285,g639,g8063,g1684,g11041,g1639,g8448,g1791,
    g8080,g248,g7323,g1707,g4907,g1759,g5668,g351,g11507,g1604,g7364,g1098,
    g6812,g932,g8570,g126,g5642,g1896,g8282,g736,g8435,g1019,g7807,g1362,g7305,
    g745,g2639,g1419,g7332,g58,g7779,g32,g11397,g876,g1086,g6808,g1486,g8444,
    g1730,g10881,g1504,g7328,g1470,g8440,g822,g8437,g583,g6291,g1678,g11039,
    g174,g8423,g1766,g7810,g1801,g8450,g186,g7317,g959,g11403,g1169,g6314,
    g1007,g7806,g1407,g8993,g1059,g7794,g1868,g7817,g758,g6797,g1718,g6337,
    g396,g11265,g1015,g7808,g38,g10872,g632,g5655,g1415,g7335,g1227,g8278,
    g1721,g10878,g882,g883,g16,g4906,g284,g7767,g426,g11256,g219,g7310,g1216,
    g1360,g806,g7289,g1428,g8992,g579,g6287,g1564,g7351,g1741,g5662,g225,g7309,
    g281,g7766,g1308,g11627,g611,g9930,g631,g5654,g1217,g9823,g1589,g7359,
    g1466,g8439,g1571,g7353,g1861,g7815,g1365,g7307,g1448,g11594,g1711,g6335,
    g1133,g6309,g1333,g11635,g153,g8426,g962,g11404,g766,g6799,g588,g6296,g486,
    g11331,g471,g11469,g1397,g7322,g580,g6288,g1950,g8288,g756,g755,g635,g5656,
    g1101,g6814,g549,g11044,g1041,g7788,g105,g11180,g1669,g11036,g1368,g7308,
    g1531,g7340,g1458,g7327,g572,g10877,g1011,g7805,g33,g10867,g1411,g7331,
    g1074,g6813,g444,g11259,g1474,g8441,g1080,g6806,g1713,g6336,g333,g5651,
    g269,g7762,g401,g11266,g1857,g11409,g9,g7336,g664,g8782,g965,g11405,g1400,
    g7324,g309,g5652,g814,g8077,g231,g7319,g557,g11048,g586,g6294,g869,g875,
    g1383,g7316,g158,g8425,g627,g5657,g1023,g7799,g259,g7755,g1361,g1206,g1327,
    g11633,g654,g8067,g293,g7770,g1346,g11656,g1633,g8873,g1753,g5666,g1508,
    g7329,g1240,g7297,g538,g11326,g416,g11269,g542,g11325,g1681,g11040,g374,
    g11440,g563,g11050,g1914,g8284,g530,g11328,g575,g11052,g1936,g9355,g55,
    g7778,g1117,g6299,g1317,g1356,g357,g11509,g386,g11263,g1601,g7363,g553,
    g11046,g166,g7747,g501,g11334,g262,g7758,g1840,g8694,g70,g7783,g318,g5646,
    g6818,g794,g6800,g36,g10870,g302,g7773,g342,g11513,g1250,g7299,g1163,g6301,
    g1810,g2044,g1032,g7800,g1432,g8990,g1053,g7792,g1453,g7326,g363,g11511,
    g330,g5650,g1157,g6303,g1357,g6330,g35,g10869,g928,g8569,g261,g7757,g516,
    g11337,g254,g7759,g778,g8076,g861,g4190,g1627,g8871,g1292,g7293,g290,g7769,
    g1850,g5671,g770,g7288,g1583,g7357,g466,g11468,g1561,g7350,g1527,g4899,
    g1546,g7345,g287,g7768,g560,g11049,g617,g8780,g17,g4894,g336,g11653,g456,
    g11466,g305,g5643,g345,g11642,g8,g2613,g1771,g7811,g865,g8275,g255,g7751,
    g1945,g9356,g1738,g5661,g1478,g8442,g1035,g7787,g1959,g4217,g1690,g6844,
    g1482,g8443,g1110,g6817,g296,g7771,g1663,g11034,g700,g8431,g1762,g5669,
    g360,g11510,g192,g6837,g1657,g10875,g722,g9346,g61,g7780,g566,g11051,g1394,
    g7809,g1089,g6809,g4897,g1071,g6804,g986,g11473,g971,g11470,g6338,g143,
    g7746,g1814,g9825,g1038,g7797,g1212,g1918,g9353,g782,g8273,g1822,g9826,
    g237,g7306,g746,g2638,g1062,g7795,g1462,g8438,g178,g7748,g366,g11512,g837,
    g4184,g599,g9819,g1854,g11408,g944,g11398,g1941,g8287,g170,g8422,g1520,
    g7334,g686,g9342,g953,g11401,g1958,g6339,g40,g10775,g1765,g3329,g1733,
    g10882,g1270,g7303,g1610,g6845,g1796,g8280,g1324,g11632,g1540,g7343,g1377,
    g7312,g4898,g491,g11332,g1849,g5670,g213,g7313,g1781,g7813,g1900,g9351,
    g1245,g7298,g108,g11593,g630,g7287,g148,g8427,g833,g4183,g1923,g8285,g936,
    g8571,g1215,g6315,g1314,g11629,g849,g4187,g1336,g11654,g272,g7763,g1806,
    g8573,g826,g8568,g1065,g7796,g1887,g8281,g37,g10871,g968,g11406,g1845,
    g5673,g1137,g6310,g1891,g9350,g1255,g7300,g257,g7753,g874,g9821,g591,g9818,
    g731,g9347,g636,g8781,g1218,g8276,g605,g9820,g79,g7776,g182,g7749,g950,
    g11400,g1129,g6308,g857,g4189,g448,g11258,g1828,g9827,g1727,g10880,g1592,
    g7360,g1703,g6843,g1932,g8286,g1624,g8870,g26,g4885,g1068,g6803,g578,g6286,
    g440,g11260,g476,g11338,g119,g7745,g668,g9340,g139,g8418,g1149,g6305,g34,
    g10868,g1848,g7366,g263,g7760,g818,g8274,g1747,g5664,g802,g6802,g275,g7764,
    g1524,g7338,g1577,g7355,g810,g7786,g391,g11264,g658,g9339,g1386,g7318,g253,
    g7750,g9822,g1125,g6307,g201,g7304,g1280,g7295,g1083,g6807,g650,g8066,
    g1636,g8874,g853,g4188,g421,g11270,g762,g6798,g956,g11402,g378,g11441,
    g1756,g5667,g589,g6297,g841,g4185,g1027,g7798,g1003,g7803,g1403,g8991,
    g1145,g6312,g1107,g6816,g1223,g8277,g406,g11267,g1811,g11185,g1642,g11183,
    g1047,g7790,g1654,g10874,g197,g6835,g1595,g7361,g1537,g7342,g727,g8434,
    g999,g7804,g798,g6801,g481,g11324,g754,g4895,g1330,g11634,g845,g4186,g790,
    g8567,g1512,g8449,g114,g1490,g8445,g1166,g6300,g1056,g7793,g348,g11506,
    g868,g1260,g7301,g260,g7756,g131,g8420,g7,g2731,g258,g7754,g521,g11330,
    g1318,g11630,g1872,g9348,g677,g9341,g582,g6290,g1393,g7320,g1549,g7346,
    g947,g11399,g1834,g9895,g1598,g7362,g1121,g6306,g1321,g11631,g506,g11335,
    g546,g11043,g1909,g9352,g6298,g1552,g7347,g584,g6292,g1687,g11042,g1586,
    g7358,g324,g5648,g1141,g6311,g1570,g4900,g1341,g11655,g1710,g4901,g1645,
    g11184,g115,g7321,g135,g8419,g525,g11329,g581,g6289,g1607,g7365,g321,g5647,
    g67,g7782,g1275,g11443,g1311,g11628,g1615,g8868,g382,g11442,g1374,g6825,
    g266,g7761,g1284,g7294,g1380,g7314,g673,g8428,g1853,g5672,g162,g8424,g411,
    g11268,g431,g11262,g1905,g8283,g1515,g7333,g1630,g8872,g49,g7774,g991,
    g7802,g1300,g7291,g339,g11505,g256,g7752,g1750,g5665,g585,g6293,g1440,
    g8988,g1666,g11035,g1528,g7339,g1351,g11657,g1648,g11181,g127,g8421,g1618,
    g11611,g1235,g7296,g299,g7772,g435,g11261,g64,g7781,g1555,g7348,g995,g7801,
    g1621,g8869,g1113,g6313,g643,g8064,g1494,g8446,g1567,g7352,g691,g8430,g534,
    g11327,g1776,g7812,g569,g10876,g1160,g6302,g9824,g1050,g7791,g1,g8078,g511,
    g11336,g1724,g10879,g12,g7337,g1878,g8695,g73,g7784,I8854,g4500,I9117,
    I12913,g7845,g11354,I17179,I10891,I10941,g6555,I6979,g2888,g5843,I9458,
    g2771,I5854,g3537,g3164,g6062,I9699,I9984,g5529,I14382,g8886,g7706,I12335,
    I13618,g8345,I15181,g9968,g6620,I10573,I12436,g7659,g5193,g4682,g6462,
    I10394,g8925,I14252,I14519,g9106,g10289,I15691,I14176,g8784,I14185,g8790,
    I16944,I14675,g9263,g2299,I12607,g7633,g3272,g2450,g2547,g9291,g8892,I6001,
    g2548,I7048,g2807,g10309,I15733,g7029,I11180,g4440,g4130,I9544,g5024,
    g10288,I15688,I12274,g7110,I9483,g5050,I12526,I6676,g2759,I8520,g4338,
    g10571,I16236,I17692,g11596,I17761,g11652,I13469,g8147,I14537,g7956,g7432,
    g3417,I6624,g4323,I11286,g6551,I8031,g3540,g7675,I12300,g8320,I13344,
    I12565,g7388,I16644,g10865,I11306,g6731,g1981,I7333,g3729,I13039,g8054,
    g3982,g3052,g6249,I10006,g9259,I15190,g9974,g11426,I17331,I14958,I13203,
    I5050,I5641,g5121,g1997,g3629,g3228,g3328,I6501,I12641,g7709,I9171,I10898,
    g8617,g8465,I15520,g10035,I7396,g4102,I7803,g3820,g3330,I6507,g2991,I6233,
    I9461,g4940,g2244,I5251,g6192,I9923,I10153,g6085,I9734,I12153,g6874,g4351,
    I7630,I11677,g7056,g10687,I16356,g4530,I7935,g8516,I13717,g5232,g4640,
    I13975,g8588,g2078,I8911,g4565,g2340,g7684,g7148,I12409,g7501,I12400,
    g11546,g11519,I10729,g5935,g5253,g4346,I11662,I7509,g3566,I9427,g4963,
    g3800,g3292,I15088,g9832,g2907,I6074,I12538,I11143,g6446,g6854,I10920,
    g11088,I16871,I11575,g8299,I13255,I9046,g4736,g6941,g6503,g2435,I14439,
    g8969,g4010,g3144,g2082,I6932,g2850,I7662,g3336,I9446,g5052,g5519,g4811,
    g5740,I9302,I5289,I9514,g5094,I12589,g2482,I5565,I5658,I15497,g10119,g2629,
    I14242,I11169,g6481,g3213,I6388,I6068,g2227,g11497,I17510,I13791,g8518,
    I16867,g10913,I10349,g6215,g10260,g10125,I12442,I8473,g4577,I14349,g8958,
    g6708,I10689,g10668,g10563,I5271,I9191,g5546,I9391,g5013,g6219,g5426,
    I15250,g9980,I17100,g11221,I14906,g9508,I14976,g7201,I11427,I14083,g8747,
    g10195,I15559,I8324,g4794,g6031,I9642,g2915,I6094,I13666,g8292,I9695,g5212,
    I11363,g6595,I11217,g6529,g6431,g6145,g6252,I10015,I10846,I14394,g4372,
    I7677,g7049,I11228,I6576,g2617,g10525,g10499,g10488,I16101,I10566,g5904,
    I13478,g8191,g5586,I8996,g8709,g8674,g2214,I9536,g5008,g6176,I9905,g4618,
    g3829,I15296,g9995,g4143,I7291,I7381,g4078,I9159,g5033,g11339,I17142,g8140,
    I13017,I16979,I16496,g10707,I12936,I7847,g3435,I9359,g5576,I13400,g2110,
    I5002,I15338,g10013,g6405,g6133,g8478,I13678,I16111,g10385,g4282,g4013,
    g11644,I17736,g7604,I12162,g9768,g9432,g4566,g3753,g7098,I11333,g10893,
    I16641,I4961,g4988,I8358,I10117,g8959,I14326,I13580,g8338,I9016,g4722,
    I6398,g2335,g8517,I13720,g3348,g2733,I15060,g9696,I15968,g10408,I5332,
    g8482,g8329,g2002,I10138,g5677,g11060,g10937,I17407,g11417,I12303,g7242,
    I9096,I15855,g10336,g2824,I5932,g11197,g11112,g4555,I7964,g5691,g5236,
    g5229,g7539,I11953,g7896,I12678,g8656,I13941,g9887,I15068,I8199,g6974,
    g6365,I10069,I14415,g8940,g3260,I6428,g11411,I17274,I10852,g6751,g10042,
    I15253,g10255,g10139,g6073,I9712,g10189,I15545,I4903,g2877,I6025,I11531,
    g7126,g10679,g10584,g6796,I8900,g4560,I16735,g10855,g1968,g5879,I9498,
    I10963,g6793,g10270,g10156,g3463,g3256,g7268,I11505,I11734,I11740,g7030,
    g10188,I15542,I12174,g6939,I12796,g7543,I9138,g7419,g7206,I15503,g10044,
    I17441,g11445,g6980,I11127,I17206,g11323,g4113,I7255,g6069,I9706,g11503,
    I17528,g7052,I11235,g8110,g7996,g2556,g4313,g3586,I16196,g10496,I7817,
    g3399,g8310,I13314,g10460,I15971,g2222,g6907,I13373,g8226,I6818,g2758,
    I7423,I6867,g2949,I9880,g5405,g10093,I15326,I10484,g6155,g9845,g9679,g3720,
    I6888,g10267,g10130,g10294,I15704,I11800,g7246,g4908,g4396,g5111,I8499,
    g11450,I13800,g8500,g5275,g4371,I11417,g6638,I17758,g11647,g3318,g2245,
    g11315,I17108,g4094,g2744,I17435,g11454,g10065,I15293,I5092,g8002,I12832,
    g5615,I9043,g4567,g3374,I8259,g4590,g11202,g7728,I12369,I10120,I14312,
    g8814,I9612,g5149,I16595,I9243,g5245,g11055,g10950,g3393,g9807,g9490,
    g11111,g10974,g4776,I9935,g5477,g4593,I8004,I11964,g6910,I7441,g3473,
    I15986,g10417,g3971,I7104,g7070,I11289,g2237,g6399,I10305,g5284,g4376,
    I11423,g6488,g7470,g6927,I15741,g7897,g7712,g7025,g6400,I6370,g2356,g7425,
    g7214,I11587,g6828,g2844,I5966,I12553,g7676,I12862,g7638,I8215,g3981,
    I10813,g6397,g11384,I17209,I14799,g9661,I6821,g3015,g2194,g10160,I15476,
    I10801,g11067,I14531,I12326,g8928,I14257,g3121,g2462,I16280,g10537,g4160,
    I7303,g3321,I6484,g2089,I4917,g4933,I8298,I14973,g9733,I5789,I16688,g10800,
    I11543,g6881,g5420,g4300,I15801,g10282,I12948,g8019,I15956,I12910,g4521,
    I14805,g9360,I10132,g2557,g4050,I7163,I13117,g7904,I12904,g7985,I4873,
    g8785,I14090,g4450,g3914,g5794,I9394,g9097,g2071,g7678,I12307,g6144,I9857,
    I11569,g6821,g3253,I6417,I7743,g3762,g6344,I10251,g3938,I11641,I15196,
    I14567,g10201,g10175,g7406,I11786,g10277,I15675,g2242,I5245,I9213,g4944,
    g3909,g2920,I6106,g2116,g7635,I12245,I4869,I13568,g8343,I13747,I15526,
    g10051,I13782,g10075,I15302,g4724,I10036,I7354,I12463,I5722,g2075,g7682,
    I13242,g8267,I17500,g11478,g6694,I10663,g4379,g3698,g3519,I12568,I11563,
    I7411,g4140,g8295,I13239,g2955,I6156,I8136,g4144,g5628,I9062,I6061,g2246,
    I12183,g7007,g6852,I10914,I11814,g7196,g5515,g4429,I6461,g2261,g5630,I9068,
    I12397,g7284,g2254,g2814,I5916,I17249,g4289,g4777,g3992,I11807,g11457,
    I17424,I9090,g5567,g4835,I8192,I14400,g8891,g2350,I5424,I12430,g9267,g9312,
    I14509,I13639,g8321,g2038,I8943,g4585,I16763,g10890,I12933,g7899,g7226,
    I11464,g8089,g7934,g10352,I15820,g2438,I11293,g6516,I13230,g8244,g2773,
    I5858,g4271,I6904,g2820,I12508,g7731,I11638,g6948,I12634,g7727,g10155,
    I15461,I17613,g11550,g10822,I16534,I4786,I6046,g2218,I9056,g4753,g6951,
    I11097,g10266,g10129,I8228,g4468,I14005,g8631,g10170,g10118,I8465,g4807,
    I16660,g10793,g7045,g6435,I10538,g5910,I8934,I5795,g7445,I11845,g6114,
    I9795,I5737,g2100,I6403,g2337,I5809,I10201,I7713,g3750,g9761,g9454,I11841,
    I11992,g7058,I11391,g6387,I9851,g2212,I13391,g8178,g6870,I10952,g4674,
    I8050,g8948,I14299,g3141,g2563,I6391,g2478,I5672,g10207,g5040,I8421,I5077,
    g1983,I10873,g3710,g3215,g7369,g7273,g7602,I12156,g10167,g10194,g10062,
    g10589,I16252,I16550,g10726,g4541,I7946,I11146,I17371,g11410,I17234,g11353,
    g7920,g7516,I11578,g6824,I12574,g7522,g10524,g10458,g2229,I15157,g9931,
    I16307,g4332,I12205,g6993,I12466,I6159,g2123,g11157,g4680,g6136,I9845,
    g8150,I7444,g4353,I7636,I10231,g8350,I13430,I13586,g8356,I15365,I8337,
    g4352,I13612,g6594,I10560,g11066,g4802,g3337,I13442,g8182,g8009,I12849,
    I5304,I15362,I6016,g2201,I6757,g2732,I12544,I9279,g5314,I9105,I10828,g5875,
    g5361,g6943,I11079,I16269,g10558,I9720,g5248,I12592,g10616,I16289,g4558,
    g3880,I9126,I13615,g8333,g7415,I11797,g7227,I11467,I9872,g5557,g10313,
    I5926,g2172,g8358,I9652,I5754,g2304,I10991,g6759,I15763,g10244,I11275,
    g6502,g10276,I15672,I17552,I8268,I7760,g3768,I16670,g10797,I11746,g6857,
    g8241,g10305,I15725,g10254,g10196,g4511,g10900,I16656,g9576,I14713,g2837,
    g2130,g10466,I15989,g5884,I9505,I5044,g6433,g5839,I9452,g8229,g7826,I6654,
    g2952,g2620,g1998,I12846,g7685,I5555,I14552,I8815,g4471,g10101,I15335,
    g10177,I15523,I16667,g10780,I13806,I7220,I5862,g2537,I9598,g5120,I7779,
    g3774,I17724,g11625,I10907,g7502,I11882,I8154,g3636,I10584,g5864,I17359,
    g11372,g3545,I6733,I15314,g10007,I17591,I15287,g6195,g3331,g6137,I9848,
    I9162,g6395,I10293,g3380,g5143,I10234,I16487,g10771,g6913,I11021,g10064,
    I15290,g11287,g11207,I15085,g9720,g2249,I9625,g4580,I10759,g5803,g11307,
    I17092,g11076,I16843,I9232,g7188,I11408,g7689,I12322,I17121,g11231,g11580,
    I11773,I10114,g5768,I9253,I9938,g5478,I16592,g11054,I10831,I9813,g5241,
    g2344,g5693,I9224,g11243,I17344,g11369,g3507,g3307,g4262,g2298,I5336,g2085,
    I7665,g3732,g10630,I16311,g11431,g6859,I10937,g7028,g6407,I6982,g2889,
    I10057,I15269,g9993,g10166,I15494,I11183,I12583,g7546,I9519,g4998,g7430,
    g7221,I15341,g10019,I5414,I16286,g10540,I7999,g4114,g2854,I5986,I17173,
    g11293,I5946,g2176,I10849,g6734,g11341,I17146,I7633,g3474,g4889,I8240,
    g2941,I6118,g6248,I10003,I17767,g9258,g3905,g10892,I16638,I14955,I14561,
    g3262,I8293,g4779,I10398,g5820,I13475,g8173,I16941,I12627,g3628,g3111,
    I10024,I7342,g6081,g4977,I10855,I10141,g5683,g4375,g3638,I10804,g6388,
    I5513,g3630,I6789,g8788,I14097,I11222,g6533,I12282,g7113,I16601,g10806,
    g5113,I8503,g6692,I10659,I16187,g10492,g6097,I9754,I7732,g3758,g7910,g7460,
    I12357,g7147,g2219,g9893,I15082,g2640,g1984,g6154,I9875,g4285,g3688,g6354,
    g5867,g2031,g10907,I16673,g5202,g6960,I11112,I15694,g10234,I5378,g2431,
    I5510,I15965,g10405,g2252,g2812,g2158,I7240,g7609,I12177,I10135,I11572,
    g8192,g2958,I6163,g8085,g7932,g10074,I15299,I8462,I13347,g8122,g9026,g8485,
    g8341,I7369,g5494,g4412,I6941,g2005,g7883,I7043,g2908,g4384,I7707,I9141,
    g5402,I9860,I8982,g4339,I9341,g10238,g10191,I16169,g10448,I9525,g5001,
    I14361,g8951,g2829,I5943,g11619,I17675,g2765,g2184,I14964,g11502,I17525,
    I12439,g2217,I13236,g8245,g7066,g7589,I12099,g4424,g3040,g2135,g4737,g3440,
    I11351,g6698,I13952,g8451,g5593,I9013,g6112,I9789,I13351,g8214,g6218,I9965,
    I10060,g3041,I10195,g11618,I17672,g9984,I15184,I11821,g7205,g10176,g10185,
    g10040,g10675,g10574,I16479,g10767,g10092,I15323,I10048,g5734,I16363,
    g10599,I16217,g10501,g3323,g2157,I15278,g10033,g7571,I12035,I11743,g4077,
    I7202,g6001,g7048,I11225,g10154,I15458,g2270,I5311,I5798,I17240,g11395,
    g7711,I12344,g4523,g3546,I10221,g6117,I11790,g8520,I13729,I17444,g8219,
    g2225,I5210,g8640,g8512,g10935,g10827,I5731,g2073,I4879,g2796,g2276,I16778,
    I6851,g2937,I7432,I7697,g3743,I10613,g6000,I11873,g6863,g10883,g10809,
    I17755,g11646,I11647,I7210,g2798,I12487,g5521,g3528,I14323,I16580,g10826,
    I17770,g11649,I16775,I8429,g2124,g3351,I6535,g5641,I9084,I17563,g11492,
    g2980,g6727,g5997,g8376,I5632,I5095,I6260,g2025,g2069,I9111,g5596,I11420,
    g4551,g3946,I15601,g10173,I9311,g4915,I15187,I12248,I13209,g8198,g4499,
    I8848,g4490,g2540,I5655,g7538,I11950,I13834,g8488,I5579,I12505,g5724,I9268,
    g9027,I14418,g2206,I5171,I12779,g7608,g10729,g6703,I10678,I9174,g4903,
    I5719,g2072,g10577,g10526,g11648,g7509,I11889,g9427,g9079,I10033,I7820,
    g3811,g4754,I16531,g10720,g10439,g10334,g6398,I12081,g6934,g5878,g5309,
    I11058,g7662,I12279,g4273,I16178,g10490,I12786,g7622,I17633,g11578,I9135,
    g5777,I9365,I10795,g6123,I13726,g8375,g7467,g1990,g2248,g8225,I17191,
    I17719,g11623,I11614,g6838,g8610,g8483,I6367,g2045,I9180,g4905,I12647,
    I16676,g10798,I16685,g10785,I11436,I9380,g10349,I15811,I14540,I16953,
    g11082,I13436,g8187,I9591,g5095,I16373,g10593,g4444,I7800,g8473,I13669,
    g2199,I17271,g2399,g9763,g7093,I11326,I12999,g7844,g3372,I10514,I12380,
    g7204,g10906,I15479,g10091,I13320,g8096,g10083,I15311,I9020,g4773,g8124,
    g8011,g10284,g7256,I11489,I12613,g8324,I13354,g11479,I17470,I6193,g2155,
    I11593,g6830,g3143,I6363,g11363,I17188,g3343,g2779,I11122,g6450,g2797,
    g2524,I13122,g7966,I6549,g2838,g4543,I10421,g5826,g6443,I6738,I6971,g2882,
    g6716,g5949,I14421,g8944,I5254,g6149,I9866,g3988,I6686,g6349,I10258,g7847,
    I12638,g3693,I11034,g6629,I10012,g5543,g3334,I6517,I5725,g2079,g7197,I9617,
    I15580,I13797,I6598,g2623,g7021,I11162,g4729,g4961,I8333,g7421,I15415,
    I5410,I8211,g5300,I10302,I10541,I6121,g2121,g1963,g110,I17324,g11347,g7263,
    I11498,I14473,g8921,g2207,I5174,g10138,I15412,I17701,g11617,I10789,I12448,
    g7530,I13409,g8141,I17534,g11495,g3792,I7017,g5353,I8820,g8849,g8745,g2259,
    I5292,g6241,I9992,g2819,g2159,I11635,g6947,I10724,g6096,g11084,I16863,
    g4414,I7752,I10325,g6003,g11110,g3621,I6754,I6938,I7668,g3733,g2852,I5982,
    I7840,g3431,I16543,g10747,g10852,g10740,I14080,I8614,g6733,I10535,I12026,
    g7119,I10434,I16938,g2701,g2040,g3113,I6343,g7562,g6984,I14358,g8950,I7390,
    g4087,I10946,g6548,g8797,I14116,g6644,I10601,g4513,g7631,I12235,g7723,
    I12354,g6119,I9810,I9973,g5502,I12616,g5901,I4920,g8291,I13227,g11373,
    I17198,g3094,I6302,I7351,g4436,I10864,g4679,I17764,g4378,g7605,I12165,
    g5511,g6823,g3518,I10682,g6051,g10576,I9040,g8144,I13027,g8344,I13412,
    g6717,I10706,I9440,g5078,I17302,I13711,g8342,I16814,g10910,I12433,g7657,
    g4335,I7612,I9123,g4890,I11109,g6464,I12418,I7363,I9323,g5620,I13109,g7981,
    g4288,I11537,g7144,g4382,I16772,g10887,g3776,g2579,g6893,g5574,g10200,
    g10169,g2825,I5935,g2650,g2006,g10608,I16283,g10115,I15353,g6386,I10282,
    g7585,I17447,I5684,I8061,g3381,g4805,g2643,I5963,g2179,I7810,g3799,g7041,
    g6427,g4005,g10863,g2008,I13606,g8311,I12971,g8039,I11303,g6526,I10081,
    g3663,g6426,I10340,g11423,g2336,I16416,g10664,g7189,g5278,I7453,g3708,
    g6170,I14506,g8923,g7673,I12296,I9655,g5173,g6125,I9822,I5707,g2418,I14228,
    g3521,I14306,I16510,g10712,g5262,g3050,I11091,g6657,g10973,I16720,g5736,
    I9296,g6382,I10099,I11071,g7669,I12286,I17246,g11543,g3996,g10184,g10039,
    I12412,g7520,I8403,g4264,g10674,g8314,I13326,g5623,I9053,I12481,I7157,
    I11255,I12133,I5957,g2178,I7357,g2122,g2228,g7531,I11929,g4095,I7233,g9554,
    I14697,I14182,g2322,I10927,g6755,g7458,g7123,g5889,I12229,I6962,g2791,
    g4495,I7886,I9839,g5226,g2230,g4437,g3345,I7244,g11514,g7890,g7479,g8650,
    I13933,I13840,I16586,g10850,g3379,I15568,g10094,g10934,g6106,I9773,g5175,
    I10177,g7505,g3878,g11242,I5098,g8008,I10240,g5937,g7011,g4719,g10692,
    I9114,I6587,I10648,g6030,I15814,g10202,g8336,I13388,I14903,g9507,I5833,
    g2103,g6121,g5285,g4355,g6461,I10391,I15807,I15974,g10411,I8858,g4506,
    g2550,g7074,I11299,g10854,g3271,I6443,g10400,g10348,g2845,g2168,I9282,
    g5633,I15639,g10179,I10563,g6043,I5584,g10214,I15586,g9324,I14970,g2195,
    g4265,g3664,g10001,I9988,g5526,I10343,g7697,g2395,g2891,I6055,g5184,I5395,
    I11483,g6567,g2913,I6088,g10329,I15775,g10186,g4442,I6985,g2890,g6904,
    I11008,g6200,g11638,g10539,I16184,g4786,g6046,I9669,I7022,I8315,g4788,
    I8811,g4465,I10370,I12981,I7118,g8289,g9529,I14672,g4164,I7311,g10538,
    I16181,g4233,g5424,I8865,I14549,g6660,I13949,g6403,g6128,g8203,I9804,g5417,
    g2859,I5995,g3997,I7131,I15510,I14570,I9792,g5403,I6832,g2909,g4454,g8033,
    I12875,I17549,g6191,g5446,g7569,I12029,I9177,g4296,I7559,I11904,g6902,
    I10633,g6015,g6735,g5231,I17318,g11340,g3332,I6513,I11252,g6542,g10241,
    g10192,g9260,g6695,I10666,I10719,I13621,g8315,g3353,I7735,g3759,g2808,
    I14191,g8795,I12953,I17616,g2342,I5406,I7782,g3775,g6107,I9776,I17540,
    g11498,I12857,g11014,I10180,g3744,g6536,I10456,I4883,g5205,g4366,g10159,
    I8880,g4537,g2255,I5276,I5728,g2084,g7688,I12793,g7619,g2481,I9202,g8195,
    g7976,I12776,g8137,I13010,I14239,g8337,g10235,g4012,I7154,g6507,I16193,
    g10485,I17377,g2097,I4935,I12765,g10683,g10612,g5742,I9308,g2726,g2021,
    I7746,I11397,g6713,I13397,g8138,g2154,I5067,g6016,I9632,I12690,g7555,I7384,
    I5070,g2960,I6173,I10861,g5980,I9567,g5556,g8807,I14140,I14573,g9029,I8237,
    I11367,g8505,g11412,I11626,I10045,g5727,g6115,I9798,g6251,I7330,I10204,
    I10843,I15275,g9994,I7674,I14045,g8603,I17739,g11641,g4787,g3423,g4728,
    I16784,I16616,g5754,I9332,g5800,I16475,g10765,g6447,g6166,I10388,g5830,
    I8234,g4232,I12445,I14388,g8924,I8328,g4801,g11305,g10972,g3092,g2181,
    I14701,g6126,I14534,g9290,g4281,g5493,g5613,g4840,I10958,g8142,I13023,
    g2112,I13406,I15983,g10414,g2267,I17698,g11616,I16766,g8255,g7986,g8081,
    g8000,g8481,g2001,g7924,g7220,I11456,g5572,I8989,g5862,I9479,I12502,I4780,
    I6040,g2216,g10522,I15517,I13574,g8360,g2329,I5383,g8354,g8717,g7023,
    I11166,I7952,g10206,g10178,I5801,I7276,g2861,g9670,I16781,g4791,I8161,
    g7977,g2828,I5940,I10075,g10535,I6432,g2727,g2022,g3736,I6924,g5534,g4545,
    g5729,I11731,g10114,I15350,I16175,g9813,I14948,I15193,g6417,I13051,g8060,
    g9987,g6935,I11065,g11193,g7051,I11232,g10107,I11756,g7191,g2221,I5198,
    g3076,I6282,I13592,g8362,g8783,g8746,g10058,I11629,I12232,g7072,I6528,
    g3274,I16264,g10557,I16790,I8490,g4526,I7420,I6648,g2635,g8218,I9658,g5150,
    g8312,I7546,g4105,I9829,g5885,g10345,g7999,I12825,g7146,I5445,I11686,
    I10162,g5943,I12239,g4049,g3375,I6569,g8001,I12829,I12261,g7078,g4449,
    g3722,I6894,I8456,g4472,g7103,I11338,g5903,g4575,g10848,I16546,g11475,
    I17466,g8293,I13233,g8129,g8015,I6010,g2256,g2068,I4866,I11152,g6469,
    I13367,g10141,I15421,g7696,g10804,I16514,I10810,g4098,g3500,I6690,I15437,
    g10050,I16209,g10452,I8851,g4498,g8828,g8744,g11437,I17362,g2677,g2034,
    g10263,g10127,I12424,I9981,g5514,g8727,g8592,g5679,I9194,g7508,g6950,g3384,
    g10332,I15782,g6213,I13837,g7944,g7410,I15347,g10135,I15403,g7521,I17164,
    I8253,I7906,g3907,g2349,I5421,g7043,I11214,I12499,g7725,I11405,g6627,g5288,
    g4438,I14528,g3424,g2896,I9132,g4893,g10361,g10268,g3737,g2834,g7443,g4935,
    g9525,g9257,I9153,g5027,I9680,g5194,I10147,g5697,I10355,g7116,g5805,I9409,
    g5916,I9550,I11596,g2198,g2231,g4268,I7523,I7771,g3418,I16607,g10787,g2855,
    I5989,g4362,I7651,g6901,I14355,I12989,g8043,g11351,I17170,g3077,g2213,
    g5422,g4470,g7034,I11191,I10825,g6588,g4419,I7763,I9744,g5263,I12056,g6929,
    g5857,I9893,g8624,g8486,g3523,g2971,I14370,g8954,g8953,I10858,g6688,I13020,
    g8049,I13583,g4452,g3365,I8872,g4529,I15063,g9699,g2241,I11394,g6056,g5947,
    I9585,I11689,g11063,I11046,g6635,I10996,g6786,I12271,g7218,g7681,g6649,
    I10610,g4746,g8677,I13962,I10367,g6234,g5824,I9901,g7101,I14367,g8884,
    g10864,g3742,I6929,g7914,g7651,g8576,I13819,g7210,I11440,I8080,I16292,
    g10551,g2644,I10671,g4730,g8716,I17546,g11500,g8149,I13036,g10947,I16708,
    g4504,I7899,I11357,g6964,g6509,I13427,g2119,I5031,I10039,g5037,I8414,
    I13357,g8125,I12199,g7278,I7372,g3226,g9311,g11422,I17321,g7035,I13105,
    g7929,I9120,g4385,I7710,g7413,g5102,I8476,g2258,I14319,g8816,g2352,I5430,
    g2818,I5922,I7140,g2641,g6063,I12529,g2175,g2867,I6007,I16635,g10862,
    I15980,g11208,g11077,I7843,I13131,I8256,I14040,I7478,g5719,I9259,g4425,
    I12843,g7683,I16717,I15235,I5388,I7435,g3459,g7936,g11542,g11453,I17416,
    g5752,I9326,I13803,g8476,g3044,I6256,g2211,g9310,I10096,g2186,I11599,g6720,
    I10713,g4637,g6118,I9807,g3983,g3222,g11614,I17662,g7601,g5265,g11436,
    g3862,g5042,I15320,I14989,g6652,g4678,g6057,I10901,I15530,g11073,g4331,
    I7606,g3543,g3101,g2170,g2614,g1994,I12490,g7922,I12712,g2125,I5053,g8319,
    I13341,g11346,I17161,I15565,g2821,I5929,g9268,I15464,I6965,g2880,g4766,
    g7033,I10739,g5942,I7249,g8152,I13043,g10421,g10331,I16537,g10721,g4305,
    g6971,g6517,g8051,I12258,I6907,I6264,g2118,I16108,g10383,g6686,I10651,
    g10163,I15485,I14010,g7597,g5296,I11249,g6541,I5638,I14645,g9088,g2083,
    I6360,g4748,I16492,g10773,I13482,g8193,I5308,g97,I11710,g7020,I12517,I4992,
    g4755,g10541,I16190,I10698,g5856,I9816,I15409,I7002,g8186,g10473,g10380,
    g4226,I11204,g6523,g6670,I7402,g4121,I17268,I6996,g2904,I7099,I13779,g8514,
    I7236,g3219,I15635,I16982,g8599,g8546,g7995,I12817,g2790,I17265,g7079,
    I11312,I11778,g3903,I7070,g5012,I8388,g9100,I13194,I10427,g4445,I10018,
    g2061,g2187,g6938,I11068,I7336,g4373,I7680,I16796,g11016,I16172,g4491,
    I12986,g7190,I11412,g8325,g6925,g7390,g6847,I12878,g5888,I13945,I12171,
    g6885,g10121,I15371,I14373,g3436,g4369,I13212,I7556,g4080,g4602,I8011,
    I11879,I17450,g3378,I6572,g5787,I9383,I9424,g5404,I17315,g11393,g10344,
    I15798,I9737,g5258,I6065,g2200,g6552,g5733,I11716,g2046,I17707,g4920,I5827,
    g2271,g2446,g4459,I17202,g11322,g3335,I6520,g8265,g8332,g4767,I8123,I7064,
    g2984,g11575,g11561,g2003,g5281,g4428,g3382,I6580,I9077,g4765,g4535,I6611,
    g2626,I8506,g4334,g2345,g10120,I17070,g11233,g8106,g7950,g11109,g8306,
    I13290,g2763,I5847,g2191,g2391,I5478,g6586,I12919,g8003,I6799,g2750,I11932,
    g6908,g3749,I14101,I9205,g11108,g2695,g2039,g9666,I14793,I12901,g5684,
    I8275,I8311,g4415,g5639,I9080,I14127,g8768,I17384,I12595,I11737,g10134,
    I15400,I7295,I11961,g7053,I16553,g10754,g5109,I8495,g5791,g3798,I13448,
    I9099,I5080,I11824,I14490,g8885,g6141,I9854,g8622,g6570,g6860,g6475,I11238,
    g6585,I14558,I5662,g9875,I15036,I13595,g9530,g6710,I10693,g5808,g5320,
    I5418,g2858,I5992,I12598,g7628,I7194,I14376,I14385,g8890,I7426,I8985,g4733,
    g11381,g4721,g2016,g2757,I5837,I13636,g7568,g5759,g5271,I10888,g6333,I6802,
    g2751,g3632,g3095,g3037,I12835,I14888,g10515,g3437,g7692,I9273,g5091,g6045,
    I17695,g3102,I4924,g3208,I6381,g7912,g8145,I13030,I13415,g2251,g2642,g1988,
    I12159,g7243,I11719,g2047,I12532,g7594,g7984,I13114,g10927,g9884,g6158,
    I9883,g3719,I12783,g7590,g11390,I17219,I13723,g8359,g5865,I9486,I13978,
    g2275,I6901,I11149,g6468,g2874,I6022,g7519,g3752,I6947,g10782,I11433,g6424,
    I16847,g10886,I11387,g6672,g5604,I9032,I13433,g8181,g5098,g2654,g2012,
    I11620,g6840,g5498,I8919,g5230,g6587,g5827,g4388,I7719,g10491,g10903,g6748,
    I13457,g6111,I9786,I10084,I10192,I7465,g10604,g8858,g8743,g4671,g3354,
    I6028,I7776,I5646,I10546,g5914,g5896,g4430,I14546,I7438,g3461,g3364,I7009,
    g5700,I8204,g3976,I12631,g7705,g8115,g7953,g4564,g8251,I13166,I13329,
    g10025,g2017,I10111,g2243,I5248,g3186,g3770,g6239,g10794,I15536,g10111,
    g10395,g10320,g5419,g9804,I14939,g10262,g10142,g10899,g10803,g6591,I10553,
    g6411,g4394,I5101,I14194,g3532,g2234,g6853,I10917,I10126,g5682,g6038,
    I16574,g10821,g4638,g2328,I12289,g7142,I6968,g2881,g6420,I10334,g11621,
    I17681,I5057,I15551,g2542,I8973,g4488,g2330,g7735,I12384,g4308,g3863,g6471,
    I17231,g11303,I12511,g6559,g5758,I12571,g3012,I6247,I11011,g6340,I5751,
    g2296,g8595,g6931,I11055,g5728,I9276,g5486,g4395,I10296,g6242,g7026,g5730,
    g5504,g7949,g7422,I7468,I16950,g3990,g2554,g4758,g4066,I7191,I13188,g10781,
    g4589,I7996,g5185,g5881,g7627,I12223,g9094,I5041,g5198,g4466,I7833,g1992,
    g6905,I5441,g3371,g11062,g7998,I12822,g10247,g4165,g4365,I13627,g8326,
    g5425,g10389,g10307,g10926,g6685,I13959,I13379,g8133,I17543,g4711,g6100,
    I9759,g6445,I17716,I10159,g7603,g4055,g7039,I9749,g5266,g10388,I8351,g8234,
    g2902,g7439,I11833,g8128,I12993,I13364,g7850,g10534,g10098,I15332,I17456,
    g4333,I7837,g4158,g8330,I13370,g10251,g10272,g10168,g2090,g4774,I7462,
    g3721,g5415,I13096,g7925,g2166,g6750,g9264,I14477,I6424,g7702,I7405,g5678,
    I10503,g5858,I16413,g10663,g10462,I15977,g3138,I6356,g8800,I14123,I14503,
    g8920,I8410,g4283,g2056,I4859,I16691,g10788,I14579,g3109,g3791,I7014,g2456,
    g7919,g7512,g10032,I15232,g2529,g2649,g10140,I15418,g4780,I8839,g4484,
    g6040,g2348,I6077,g11574,g11452,I17413,I16802,I9199,g5766,I9346,I8487,
    g4509,g6440,g6150,g1976,g11205,I6477,g7952,g7427,g9450,g5305,g5801,I5734,
    I6523,I4820,I17243,g11396,I5435,g2851,I5979,g2833,I12559,g7477,I14315,
    g8815,I6643,g3008,g8213,I10819,g6706,g11311,I10910,I9102,I9208,g5047,g3707,
    I14910,g9532,g7616,I12196,g7561,I12015,g4067,I6958,I8278,g8805,g5748,I9320,
    I10979,g6565,g2964,g4418,I9869,g4467,I15072,g9713,I14979,g9671,g4290,
    I14055,I16583,g7004,g11072,I17773,g11650,I15592,I15756,g7527,I6742,g3326,
    g4093,g2965,I8282,g4770,g6151,I12457,g4256,g6648,I10607,g9777,g9474,I11970,
    I10384,g5842,g10162,I15482,g3715,I9265,g5085,I16787,g10896,g11350,I5713,
    g2436,g10204,g8056,g7671,I13317,g8093,I12610,I7360,g2906,g8529,I13738,
    I14094,g8700,g4381,g7476,g5396,g8348,I13424,I12255,g7203,I6273,g2872,
    I16105,g10382,g10629,g10583,I10150,g5705,g5169,g4596,I7408,g8155,I13048,
    I13002,g8045,g8355,I13445,g10220,g5007,I8379,I13057,g7843,g2652,g2057,
    g7376,I13128,g2843,g10911,I11608,g2989,g3539,g4263,I13245,g8269,g7042,
    I16769,g10894,g5718,I9256,I12460,I12939,g5767,I9349,g10233,I13323,I7176,
    I5976,g2549,g2853,I10526,g6161,I12907,I5952,g6172,I10093,g7617,g3861,g7906,
    I12694,I17258,g5261,g10591,I16258,I6543,g3362,I6546,g3419,g3104,I7829,
    g3425,g6667,I10630,g4562,I7973,g6343,I10248,I16439,I14564,g10355,I15829,
    I10105,I12478,g6566,g7027,g4631,g10825,g6732,I15583,g10157,g9802,g1999,
    g6537,g4257,g6134,I13338,I14188,g5221,g2232,I5221,g10172,I16799,g3086,
    g5203,g2253,g3728,g2813,I5913,I9029,g4781,I14077,g8758,g4902,g6080,I9371,
    g5075,I10822,I15787,g10269,I6414,g3730,I6080,I9956,g5485,g6059,g3385,
    g11357,I17182,g7991,I12809,g10319,g4441,g6113,I10198,I11309,I11668,I10102,
    g10891,I13831,g8560,g10318,I15752,g4089,I5588,g8121,I12978,g10227,g7907,
    g7664,I6436,g2351,I6679,g4673,g6202,g8670,g8551,g5689,I9216,g4757,I9684,
    I11194,I15768,g10249,g5210,I9639,g5126,g7959,I12751,I10066,g5778,I9338,
    g8625,g8487,g7082,I11315,g2586,g1972,g5216,I17410,g11419,g6094,g6578,
    I16647,g10866,I15281,g10597,g4669,I8724,I10495,g4368,I11989,g6919,I17666,
    g11603,I10885,g6332,g4231,I6510,g10203,I14876,g9526,I11611,g7656,I12265,
    g4772,g3406,I11722,I7399,I15263,g3635,I6812,g4458,g2570,g2860,I5998,g2341,
    I5403,g9262,g3682,g6593,I10557,g5344,g8519,g3105,g7915,g7473,g3305,I6474,
    g10281,g98,I4783,g2645,g1991,I8835,g7677,g10902,g8606,I11450,I15368,g4011,
    I7151,g9076,g5741,I9305,g3748,g4411,g4734,I11342,g9889,I11345,I10051,I6560,
    g3212,I8611,g5844,g5638,g6933,I11061,g7663,I11650,g10699,I16376,I12853,
    I16897,I5240,g2962,I6183,g6521,I10437,I17084,g11249,g4474,g10290,g6050,
    I9677,g6641,I10598,I11198,g5081,g10698,g2506,I10378,I6037,g2560,g11348,
    g5883,I10314,g7402,I6495,g2076,I9833,g5197,I11528,I6102,g2240,g10779,
    I17531,g11488,I7694,I11330,g6571,g3373,I6565,I15778,I12451,g3491,g2669,
    g2903,I5116,g11081,I16856,I7852,g3438,I7923,g3394,g5066,I8436,g5589,I9001,
    g6724,I13403,I10054,I9539,g5354,I9896,g5295,g4713,I10243,g5918,I11132,
    g6451,I11869,g6894,g7877,I7701,g3513,g3369,I6557,I6240,I14522,I15356,
    I12268,g6878,I10966,I15826,g10205,I6917,g2832,I15380,I4894,g2174,I6661,
    g9024,I14409,g2374,g7534,g5035,g7556,I16723,g10851,g3767,I6976,g10547,
    I16206,g9424,g10895,g4076,I9362,g2985,I6217,g9809,I14944,I9443,g6882,
    I10974,g7928,I10156,I10655,g6036,g10132,g3582,I16387,I17334,g11360,I10072,
    g6534,g10226,I15598,I16947,g11651,g7064,I11269,g2239,g9672,I13708,g5774,
    I12683,g3793,g2593,g7464,I11858,I12053,g6928,I13454,g7686,I12520,I16811,
    g10908,I16214,g3415,g3227,I6406,I7825,g3414,I10807,g2171,I11043,g6412,
    I6454,g2368,g8055,I17216,g11291,g2420,g6674,I10639,I17558,g7259,I15383,
    g3209,I13197,g2507,g3246,I15448,g10056,g5509,g4739,g4326,I14694,g4125,
    g7237,I11477,I9185,I6891,I11602,g6833,I11810,I17255,g6132,I9147,I6553,
    I4850,g11499,I13068,g6680,I10643,g6209,g5994,g10889,I16629,I16850,g10905,
    g6918,g7394,g6197,g10354,g2905,g7089,I11322,I12376,g10888,I16626,I10816,
    g8239,I7366,g9273,g4608,g3726,I12762,I4948,I10278,g5815,g3940,g6558,I12009,
    g6915,I8262,g4636,I11967,g6911,g8020,I10286,g6237,I5060,g10931,g3388,I6590,
    g8812,I11459,g11433,I17350,g9572,I14709,g5685,I9237,g8794,I14109,g5397,
    I5818,I8889,g4553,g11620,I17678,g10190,I15548,g4361,I7648,I9766,g5348,
    g3428,I6639,I7096,I12454,g7544,I9087,g4970,I9801,g5416,g3430,g7441,I17742,
    g4051,I7166,g5996,g8047,g11343,I17152,I13918,I16379,g10598,g4127,g4451,
    g4327,I7600,g11352,I11698,g6574,g2196,g10546,I16203,g7038,I11201,I11444,
    g6653,g11420,g10211,g9534,I14687,I15162,g6714,g7438,g7232,I12484,g6832,
    g7009,I17194,I5047,g2632,I7625,g8515,I13714,g10088,I15317,I8285,g4771,
    g7073,I5840,g2432,g9990,g11481,I16742,g10857,g8100,g7947,g11079,g3910,
    I13086,I12472,I8139,g3681,g7212,g5723,I14884,I17277,I11817,I10168,g5982,
    g5817,g7918,g5301,g7967,I15229,I5427,I11159,g6478,g10700,I5765,I9491,g5072,
    g10126,I8024,g4117,I11901,g6897,g2530,g6736,I13125,g7975,g8750,g6042,g4508,
    g10250,g10136,g2655,g2013,g4240,I11783,I16793,I9602,I5704,g7993,I12813,
    g6076,I9717,I4906,I11656,g7122,I6049,g5751,I6955,g3066,I8231,g4170,g4443,
    g3359,g10296,I15708,I11680,I14340,I17116,g11229,g2410,g9452,I7726,g6175,
    g4116,I7260,g6871,g2884,g2839,I7054,I6498,I17746,g11643,g3055,I15959,
    g10402,g7921,g7463,g10197,g4347,I8551,g4342,g3333,I9415,I17237,g11394,
    g4681,g4330,I12577,g7532,g8151,g8036,g10527,I6999,g8351,I17340,g11366,
    g4533,I7938,g7848,g8221,I15386,g6184,I9915,g2235,g2343,I9168,I10531,g6169,
    I17684,g11609,I14179,I7447,I7112,g11301,g11096,I16879,g7620,I12208,I8007,
    g3538,I6726,I6019,g6140,g10859,I10186,g6110,g6737,I16571,g2334,I10837,
    I10685,g6054,g5743,g4413,I7749,g5890,g6508,I6052,g2220,I5667,g8956,g6531,
    g8050,I14224,I16298,g10553,I13224,g8261,g6077,g11429,g5011,I8385,g3067,
    I13571,g10315,g10243,I9290,g10819,I16525,g11428,I17337,I16682,g3290,g11376,
    g10171,g10257,g4317,I7586,I13206,I4876,g3093,I6299,g5474,g7192,g6742,g5992,
    I9608,g7085,I11318,g3763,g6634,I10589,I9188,I10762,g6127,g8667,g3816,g8143,
    g8029,I13816,g8559,I6504,g3214,I9388,g8235,g11548,g6104,I9769,g9762,g10590,
    I16255,I6385,g2260,I10171,g10909,g6499,I16261,g10556,g2202,g11504,g4775,
    I11752,g7032,g8134,I13005,g7941,g8334,I13382,g9265,g2094,I12415,g11317,
    I17112,I15329,g3397,g8548,g8390,g2518,g4060,g4460,I9564,g3697,I10078,I8885,
    g4548,g8804,I14133,I14543,g4293,g10150,I16507,I9826,g5390,g7708,I12339,
    g8294,g10735,g11057,I11898,g8792,I14105,I17347,g3735,g6044,I9665,g1973,
    g7031,g6413,I8903,g4561,g6444,g11245,g7431,I12601,g11626,g9770,I15562,
    g6569,g10695,I16366,g5688,I17124,I13489,g8233,I6196,g2339,I5475,I7716,
    g3751,g6572,g6862,I5949,g7580,g8787,I9108,g10253,g8200,g4479,I7858,I14681,
    g6712,g5984,I8036,g4294,I10123,g5676,g6543,g4462,g9553,g8767,g3723,g3071,
    g7286,I11534,I7387,g2197,g4390,g6396,I15962,g3817,g7911,g6563,g8094,g7987,
    g2050,g1987,I8831,g4480,I17516,g11483,I16432,g10702,g4501,g6729,g6961,
    I11115,I13794,g5863,g4156,I11713,g7733,I5850,g2273,g7270,I11515,I11049,
    I6944,I9165,I16461,I9571,g5392,g7610,I12180,g4942,I8308,I14424,g6014,
    I11296,I12799,g9429,g9082,g22,I4777,g5838,g11289,I10623,g6547,g10256,
    I17555,g8270,I14391,I16650,g10776,I6373,g2024,I6091,g5183,g7124,g7980,
    g10280,g6903,I11005,g2777,I5919,I11188,g6513,g7069,I12805,g8171,g5779,
    g9272,g4954,g4250,g4163,I7308,I6034,g7540,I11956,g8160,g4363,I7654,I16528,
    g10732,I7577,g4124,I13460,g10898,g5423,I17453,g11451,I11383,g6385,g7377,
    I11759,I15467,I9647,I5561,g8052,g4453,I13648,g6178,I6767,g2914,g4325,g3368,
    g9745,g2826,g2799,I17513,g6135,I9842,I9156,g9109,I14452,I10228,g9309,g3531,
    I8869,g4421,g5127,I8535,g3458,g6182,g11389,I9662,g5319,g8179,g7849,I12644,
    I16598,g10885,g11056,g8379,I13485,g4912,g8766,g2997,I17657,g7537,g2541,
    g11080,I16853,g5146,g10708,g3505,I6694,I5970,g2185,g6749,I10756,g2238,
    I5237,g11432,g3411,I6616,I9093,g7900,g10555,g2209,I12556,I8265,g5696,I9229,
    I11085,I7984,I5224,I7280,I10237,g6120,I8442,g4464,g7658,I13185,g2802,
    g11342,I17149,g6205,I5120,g9449,g6560,g8820,g5753,I9329,I8164,I15736,
    g10258,g10456,g5508,I8929,g11199,I14684,g9124,I17752,I11617,g6839,I13915,
    g5472,I14364,I9421,g5063,g2162,g5043,g6522,g10314,I15744,I11494,g5443,
    g6208,I9953,I7790,g3782,g10936,I10165,I15729,I7061,g6579,g5116,g6869,
    I10949,g7852,g7923,g11320,g4083,g10596,g8339,g8132,g6719,I10710,I13376,
    I11623,g6841,g7387,g8680,I13965,g10431,g10328,I11037,g8353,I13439,I14130,
    g8769,I10362,g6224,g2864,g5948,g6917,I11029,I8247,g2208,g8802,I6671,g7886,
    g4735,I17327,g11349,I7109,g4782,I11155,g6470,I17537,I13418,I13822,g6442,
    I11590,I8631,g11225,I7345,I16458,g10734,I9605,g4475,g6164,g3769,g2646,
    g5755,g10335,g7650,I15244,g10031,g4292,g10930,g6454,g11244,I7931,g6515,
    g3760,g3003,g7008,I13589,g8361,I17381,I7536,I4886,g10131,I15395,I11524,
    g11069,g4084,g3119,I11836,g4603,g5936,g8600,g8475,g9710,I12469,g4439,I7793,
    g5117,g6553,I10477,g8714,g11068,g3631,I12120,g10487,I16098,g7972,I12770,
    I11119,g9025,I14412,g2871,I6013,g10619,I12759,I7757,I16817,g10912,I9673,
    g5182,I14236,g6556,g3220,I8109,g3622,g2651,g2007,g2302,g4583,I10322,I17390,
    g11430,g10279,g10158,g7065,I11272,I7315,g6389,I10289,I7642,g7887,g7693,
    I15792,I9368,g4919,I8290,I10063,g6990,g3694,g10278,g10182,g3977,I6861,
    g2942,g6888,I10984,g10791,I9531,g5004,g6171,I16295,g10552,g3161,I11704,
    g7632,g2569,I17522,g11485,I5399,g6331,g6956,I11106,g5597,I9023,I14873,
    I13809,g8480,I6133,g3051,g2165,I12930,g10069,I13466,g5088,I13674,g2424,
    I8449,g4469,I12652,g9766,g2809,I5909,g5784,g4004,g5257,g8053,g4518,g7550,
    I11560,g7037,g10187,I15539,I5824,g2502,I10834,g6715,g3633,I15079,I8098,
    g3583,g2077,I5218,g7195,g11545,g11444,g7395,I13642,g8378,I11659,g3103,
    I9074,g4764,g7913,I6538,g2827,g2523,I7272,g1989,g10143,I15427,g11078,
    I10021,g5692,g5840,I13695,g11598,I17642,g3068,g6109,I12406,g11086,I12586,
    I7417,I6914,I17252,g8184,g10884,I15817,g10199,I9863,g8139,g8025,g2742,
    g3944,I15500,g5763,g6707,I13630,I5348,g9091,g4320,g11159,I10274,g5811,
    g6480,I11665,g3761,I5064,I14112,g10217,I15589,g4277,g6201,I11674,g6795,
    g6957,g2754,I5830,g4789,g10486,I16095,I17176,I15823,g6449,g8194,g8477,
    g8317,g6575,g7525,g8523,I13732,g2257,g9767,I14914,g7097,I9688,g5201,g7726,
    I12363,g5269,g8183,I5740,g7497,g9535,I14690,I10702,g10580,g10530,g2444,
    g5032,g2269,g10223,I15595,I7213,g9261,I6421,g2346,g4299,g8938,g7579,I6856,
    g8099,g7990,g4238,I14136,g8775,g8304,I13280,g4891,g8266,g10110,I15344,
    g2543,g6584,g11017,g6539,I10461,g6896,g5568,g10321,I15759,I5089,I17213,
    g11290,I12514,g10041,g10531,g10471,g7979,g3413,g5912,I11584,g4738,I11519,
    I11176,g6501,g7001,I11140,I13191,g10676,g10570,g6419,I10331,g6334,I7456,
    g3716,g1993,I7284,g6052,g11309,I17096,I7205,g8613,g8484,g10719,I7348,g4056,
    g6452,I15308,g4478,g2014,g2885,I6043,I9779,g5391,g2946,g4435,g4727,g4082,
    I12421,g7634,I8406,g4274,g8765,I12366,g3433,g9308,I10108,g6086,g8712,
    I12012,g6916,I9588,g5114,I12403,I5438,g11377,I14303,g8811,I10971,I12541,
    g7703,g5174,g10264,I5525,I15374,g9028,g8729,g8961,I14330,I4900,I11501,
    g6581,I16610,g10792,I14802,g11308,g3060,g8290,I13577,I10381,g5847,I7459,
    g10554,I14982,g6425,I11728,g7010,I17733,I16679,g10784,I5391,g2979,g4310,
    g2382,I7318,g3266,g7680,I16124,g10396,I12535,I10174,I15669,g10543,g3784,
    g11425,g5894,g10117,I15359,g8660,g8946,I14295,g2916,I6097,g5735,I9293,
    I15392,g10104,g2749,I5815,g3995,g3937,I7086,I10840,g9741,g4002,I7393,g4096,
    I6531,I11348,g7062,I13083,g3479,g11195,I17482,g6131,g5548,I9144,g8513,
    I15488,g10116,I15424,g10080,g6406,g10242,I15632,g5475,I8892,g4762,I8116,
    g2449,I11695,g11424,I9240,g5069,I10592,I11566,g6820,I16739,g9108,I14449,
    g3390,I14499,g5627,g5292,g9883,g3501,g4340,g5998,I9620,I13385,g2873,I10753,
    g2095,I11653,g6954,g2037,I13099,g4222,g5603,g2297,g5039,I8418,I4951,g10293,
    I15701,g2653,g2011,g6922,g5850,g6226,g3704,g10265,g1969,g8357,g6747,g11391,
    g2719,g2043,g9448,I7909,g3387,g2108,g8818,g4785,g10391,I6480,g5702,g2752,
    g8649,g9555,g6091,g6071,g3810,g3363,I10904,g8798,I14119,I11354,I11605,
    g3432,g10579,g10528,g4563,g9774,g4166,I13773,I16277,g10536,g2042,g4295,
    g10578,g4237,I10317,g6868,g5616,g10783,g8632,g8095,g7942,g2164,g6718,g2364,
    g2233,g9780,I16623,g10858,I13609,I10183,g6108,g11065,I7729,I5192,g2054,
    g6582,I14397,g8888,g7386,I11767,g4731,I8085,g2454,I5549,g8579,I12773,
    I13200,I10042,I12604,g7630,g8719,g4557,I9317,g2725,g2018,g1974,g8926,
    I11173,g4239,g4966,I8340,I14933,g7426,I14494,I11921,g11602,g8041,g8752,
    g8635,g6227,g5503,g4515,g7614,I12190,g10275,g4242,g10493,I16114,g4948,
    I7691,g9816,g1980,g4615,g11160,I13624,I17710,g6203,I9581,I15241,g4254,
    I16589,g10820,I16518,g8164,g7872,I15470,I5812,I17669,g2131,I7659,g3731,
    g7636,I6220,I4891,g8922,I8133,g8296,g2956,I15075,g8725,g8589,g3683,I6844,
    g11075,g2004,g10165,g10079,I17356,g8532,I13741,g7187,g2803,g4769,g5987,
    I11692,I11770,I17438,I9995,g5536,g6689,I17687,g10193,g10057,g10796,g5299,
    g4393,g5810,g10259,g7067,I6921,I15491,g8236,g10523,g11605,I7006,I13013,
    g8048,g5892,g6528,I17312,g2745,g2338,I5073,g8116,I11207,g6524,g7446,g3475,
    g3056,g11155,g3255,I15266,g7258,I12388,g7219,g8046,I14232,g7403,g3627,
    I6784,g4822,g3706,I12871,g6564,I16808,I11683,g11482,I8711,g2156,g2373,
    I12251,g7076,g10381,g2707,g2041,I8827,g4477,g10437,g10333,I5843,g4456,
    g4167,g7637,g10161,g3039,g2310,g3439,g7107,I12032,g6923,g8297,g10347,I8396,
    g4255,g3624,I11725,g5082,g4732,I11100,g5482,I14405,g8937,g10600,g4752,
    g8684,I13969,I8250,g5876,g2363,g6538,I13394,g10236,g4062,I7185,g2098,I4938,
    I9129,g7416,g4620,g10351,I15864,g10339,g6589,I10549,g3524,I15749,g2210,
    g11306,g7047,I7300,g2883,g11313,I17104,I12360,g7183,g4778,g10063,I17387,
    g11438,g8707,g8671,g6165,g10128,g6861,g5214,g10137,g6048,g9772,g6895,g2539,
    I5652,I6347,g6448,I10374,g9531,I14678,I15305,g6711,g6055,g11223,g11053,
    g9890,g6163,g3404,I9836,I9150,g6179,g9505,g9052,g9721,g2268,I13645,g4298,
    g3764,g8575,g8776,g4485,I8842,g6196,g7880,g7595,I12123,I11947,I17368,g8604,
    g8479,g10208,I16239,I17730,g8498,g6827,g4309,g9331,g7272,g8197,g10542,
    g11064,g7612,I12186,g2086,g7244,g7040,g7586,g2728,g7930,g6418,I11082,g7982,
    I12790,g4520,g5222,I17228,g11300,I17704,g4219,I10129,I6031,g4061,g10718,
    I6601,g3727,g7629,I15665,I11632,g2070,g3906,g11622,I13744,g10346,I15804,
    g5899,g4958,I10027,g10122,I7143,g10464,g10034,I15238,g6181,I11804,I14249,
    I17419,g6482,g10292,I15698,I9475,g5445,I9930,g6700,g11227,g6088,I10299,
    g7213,I11447,g2331,I16577,I8089,g2406,I13332,g8206,g4270,I11135,g6679,
    g4057,I15406,g11636,I12318,g11074,g10901,I11094,g11239,g11219,g4225,g2087,
    I17636,g3945,g2801,g2117,g5089,g4886,g3738,g3062,I14786,g9266,I12867,g9760,
    I6294,g11608,g3709,I6870,I7269,g4324,g2748,g6562,g10164,g7077,g10133,I9248,
    g5471,g4370,g2755,I16956,I7076,g2226,g2578,I10090,g6723,I10716,g8059,
    I10030,g8771,g11518,g6101,I9762,g7649,g2459,g4377,g6035,g3517,I6702,g10575,
    g7851,g11501,g3876,g8131,g10327,I15771,g2173,g7106,g4287,g6198,g7964,
    I12562,g8105,g7992,g2169,g8973,g10283,g2369,g6834,I7414,g5773,g4399,g6921,
    g2407,I14961,g9769,g1962,g2868,I8147,g6041,g2647,I13812,g5148,g6441,I13463,
    g8156,I14642,g3110,g11577,g7279,g5836,g4510,I12427,g7134,g2793,g4291,
    I12655,I17365,g10174,I15514,I16500,I16664,g10795,g9103,g2015,g6368,I13633,
    g3773,g7057,g4344,I5142,I7593,g4142,g7989,I15284,g7611,I12547,g11083,
    g11276,g10390,I16484,g10770,g9732,g5218,g11284,g5822,g4819,g3877,g9271,
    I12226,g8007,I7264,g3252,g2203,I15554,I10620,I5497,g2846,g7570,I13421,
    I16200,g10494,I5960,g4081,g8773,g6856,I10924,I10733,g5401,g8535,I7450,
    g8582,I13825,g7670,I17261,g3462,g4951,I8320,I11472,I16220,g5895,g7938,
    I8126,g3662,g4314,g5062,I13788,g10326,g4417,g7909,g2689,I12103,I11829,
    g6740,g10484,I16805,g10904,g8664,I15247,I10412,g5821,g7143,g9533,g8939,
    I13828,g2028,g8772,g10252,g8721,I10499,g10621,g7606,I12168,g2247,I5258,
    g4336,g2067,g2564,g7687,g4768,g11576,I17610,g6093,I13682,I6911,g2163,g6500,
    g10183,g5192,g4943,g3352,g11200,g3705,g10500,g11388,g4065,g2794,g3637,
    g4228,g4322,g5941,I14379,g4934,g4243,I11671,g6485,I10308,g8777,g6244,
    I13956,I6439,g5304,g3254,g9775,g11640,g3814,g5708,g5520,g11319,I13785,
    g3038,g1982,g4496,I7889,I8303,g4784,g5252,g7607,g11487,g5812,g3009,g9110,
    g6183,g2571,g5176,g6220,I5716,I5149,g10047,g4337,g4913,g11380,g2055,g10311,
    g2455,g9739,I6952,g9269,I9402,g5107,g7054,g4380,g1975,g7236,I11581,g2774,
    g3967,g3247,g11314,g7729,g5276,I15272,g9150,I9886,g7615,I12193,g6361,g4266,
    g4159,g9668,g2396,g10592,I9287,I17225,g11298,g7202,g5270,g4367,g7374,g6819,
    I12916,g11345,I7288,g2509,I16407,g10696,g2987,g5073,g10350,g11539,g6146,
    g7545,g2662,g5124,I9594,g7380,g6103,g5317,I11794,g8711,g7591,g8472,g4726,
    g2994,g5469,g7853,g4354,I7639,g7420,g5177,g8346,g11241,g10453,g6243,I5279,
    g6514,g7559,g8817,g10691,I16360,g8810,g8196,g6944,g8803,I6277,g6072,g8538,
    g2381,g9313,g10387,g4783,I7375,g2847,I5973,g6157,I12202,g6983,g8509,g8366,
    g9453,g4112,g7905,g7450,g4312,g4473,g6577,g10929,I12496,g7724,g5195,g6116,
    g2421,g4001,g3200,g8040,g10928,I9731,g5255,g5898,g6434,I10352,g4676,g5900,
    g5790,I5821,g2101,I11926,g6900,g8042,g4129,g5797,I9399,g4329,g4761,g11515,
    g11490,I7339,g7927,g8230,g6681,I11701,g5291,g3392,g6546,g3485,g2562,g6697,
    g5144,g4592,g6914,I11024,g11446,g6210,I12150,g6596,g4221,g8381,g2817,g3941,
    g7440,g8574,I10445,g5770,I17374,I11360,g8889,g7648,g5701,g4953,g3520,
    g10711,I6395,g2743,I15114,g9719,I17158,g11312,I16613,g11435,I6876,g5287,
    I16859,g3812,g5886,g11107,g6351,g10261,I13360,g8126,I17353,g3405,g9778,
    g4387,g9894,g8723,g8585,g4716,g6479,g3765,g3120,g5814,g5849,g3911,I16632,
    g9782,I5695,I5111,g6060,I16273,g10559,g5219,g4747,I10736,g4398,I13451,
    g10248,g2772,g2508,g7240,g8751,g4241,I9352,g5594,g9270,g8819,g9256,g6656,
    g6995,g7618,g3980,g2411,I5494,g10786,I13776,g4524,g3757,g5887,I9510,g10356,
    I15832,g5122,I17519,g6190,g2074,g4319,g6906,g10717,I16540,g4759,g3206,
    g5189,g4258,g4867,g6156,g4717,g2919,I10087,g9919,g2080,I14087,g8770,g2480,
    g6392,g6621,g5096,I11076,g2713,g6704,g11610,g4386,g10932,g4582,g5845,g4975,
    I7513,g11645,g5395,g5891,g11106,g4426,g10897,g6250,I10009,g4614,g9527,
    I14668,I7671,I12550,I7378,g6432,g7908,g7454,g8264,g6053,g9765,g11604,g9764,
    I16920,I16760,g3291,g2161,g7245,g6453,g4280,I7182,g4939,I11540,g6877,g2510,
    I15795,g3344,I16121,g6568,I7216,I12942,g4544,g3207,g2439,I7916,I12493,
    g2000,g8713,g11486,g2126,I6071,I14967,g7581,g10799,I15507,g3088,g4306,
    g7965,g5481,g4790,I9221,g1964,g10357,g7264,g10620,g10148,g11421,g4461,
    g6439,g4756,I17713,g8688,g8507,g7133,g10343,g8642,I14918,g4427,g8044,
    I15473,g10087,g8254,I6150,g11541,g11549,g9771,I12838,g2023,g11344,g4514,
    g5874,g5783,I9377,g4003,I6409,g5112,g7379,I8647,g11232,g5267,g11607,g6573,
    g9892,I8039,g3506,g3407,g4763,g7878,g8760,g11434,g4391,g6193,g3408,g3108,
    g2451,g7225,g6778,g7882,I17155,g4307,g4536,g10228,I15604,g4359,I13102,
    g8608,g8220,g7231,g4576,g3943,g4904,I10144,I14525,g8806,g11292,I16604,
    g6822,g4416,g7624,I14352,I5792,g10310,g7997,g2753,g4315,g3661,I15861,g6561,
    I11644,g10378,I15858,g5624,I11707,g6084,g8327,g8952,g4874,g6039,g5068,
    g6912,g3096,I11103,g3496,g6898,g8146,I5020,g5421,g8103,g7994,g3395,g2434,
    g3913,g6583,g6702,g4880,g5866,g8696,I7029,I14309,g8813,g2347,I7429,g10802,
    I7956,g7901,g4272,g10730,g7560,g6924,I17749,g8240,g5747,g4420,g5308,g7600,
    I12580,g7574,I6085,g10548,g11310,g3142,g6527,g4328,g11294,g3815,I11211,
    g5852,g6764,g2970,g6026,I11088,g9556,g10369,g10317,g3097,g5286,I6898,g6970,
    g2317,g4554,I15389,I15127,g3370,g5818,g8697,g8024,g10323,g11191,g2775,
    g3783,g5893,g5106,g8945,g3112,g3267,g7983,g4804,g6525,g2060,g6617,g6019,
    g6789,g8210,g5083,g3585,g11573,I5710,g5614,g7541,I7173,g7500,I13335,I9433,
    g3828,g10697,I16370,I9065,g4760,g11447,g8601,g2479,g10860,g2840,I10189,
    g7024,g10502,g2190,g4260,g2390,g11579,g7737,g3703,g4463,g7672,I12293,g6709,
    g11639,g9814,g5030,g6826,I14555,g2303,g8739,I12242,g4279,g9773,g11061,
    g10498,g9009,g6082,I9727,g4318,g4872,g7626,g5200,g4457,I8877,g6829,I17185,
    g10271,g9958,g4549,g7211,g11162,g5191,g3747,g10342,g3398,g6214,g10145,
    I9783,g5637,g7044,g2912,I13735,g8704,g4321,g10198,g5223,I7487,g7660,g8363,
    g10330,g10393,I7766,g10722,g6236,g11071,g8887,g11484,g11286,g6002,g11606,
    g11217,g10454,g4519,I7920,g5251,g6590,I11942,I12372,g7961,g6757,g4552,
    g4606,g6216,g8941,g10856,g7414,g3386,g4892,g7946,g3975,g4586,g7903,g2683,
    g3426,g5880,g6930,g8250,g2778,g5250,g5272,g7036,g9085,g4525,g7436,g8626,
    g6049,g8943,g10861,g11059,g2475,g8779,g3544,g11540,I6815,g5629,g5484,g6089,
    g7916,g11203,g5542,I8967,g7022,g3306,g2998,g3304,g6557,I12523,g3790,g4482,
    g6705,g5190,g6180,I15377,g9431,g9812,g3756,g4587,I12475,g5274,g4275,g4311,
    g3427,g5213,g8774,g10545,g10444,g10325,g7437,g8260,g4284,g8526,g6099,g3391,
    g10401,g5490,I14485,g11427,g5166,g6831,g4591,g6068,g7137,g7917,g9473,
    g10532,g1965,g4507,g6967,g6545,g2764,g11547,g7257,g6909,g8384,g7442,g8702,
    g2503,g11392,g10353,g3416,g6506,g8883,g3522,g11572,g2224,g6728,g10724,
    g2320,g4556,g3070,g3874,g8004,g2789,g5619,g5167,g11103,g2250,g9900,g11095,
    g4973,g7389,g7888,g7465,g4969,g8224,g2892,g5686,g10308,g4123,g8120,g6788,
    g5598,g4824,g9694,g10495,g2945,g11190,g8789,g8639,g9852,g9728,g9563,g5625,
    g4875,g9701,g7138,g10752,g11211,g11058,g11024,g8547,g8307,g10669,g7707,
    g4884,g3813,g4839,g9870,g6640,g9650,g9240,g5687,g7957,g3512,g7449,g4235,
    g4343,g11296,g9594,g9292,g9943,g9923,g9367,g5525,g8876,g10705,g10564,g9934,
    g9913,g9624,g6225,g6324,g10686,g6540,g8663,g11581,g6206,g3989,g7730,g7260,
    g7504,g7185,I5689,I5690,g7881,g11070,g9859,g9736,g9573,g8877,g11590,g2274,
    g6199,g8932,g5545,g5180,g5591,g8556,g8412,g11094,g5853,g5044,g6245,g4360,
    g8930,g5507,g11150,g3087,g8464,g8302,g9692,g4996,g7131,g11019,g9960,g9951,
    g9536,g11196,g11018,g10595,g10550,g10433,g10623,g10544,g4878,g5204,g4838,
    g8844,g8609,g6701,g6185,g10725,g5100,g4882,g8731,g5128,g6886,g8557,g8415,
    g8966,g8071,g11597,g9828,g9722,g9785,g2918,g9830,g9725,g8955,g9592,g5123,
    g7059,g6078,g7459,g11102,g7718,g7535,g9703,g5528,g5151,g9932,g9911,g5530,
    g2760,g8629,g6887,g6187,g6228,g5605,g6322,I6337,I6338,g8967,g5010,g3275,
    g2895,g7721,g9866,g9716,g10808,g10744,g3047,g4492,g3685,g8822,g8614,g10560,
    g11456,g9848,g9724,g9557,g4714,g6550,g5172,g10642,g3284,g2531,g9855,g5618,
    g6891,g7940,g11085,g4968,g8837,g8646,g9644,g9125,g5804,g8462,g8300,I6330,
    g11156,g6342,g9867,g9717,g4871,g10435,g7741,g9386,g9151,g8842,g8607,g9599,
    g9274,g8974,g5518,g9614,g9111,g4122,g7217,g4610,g11557,g2911,g11210,g7466,
    g9939,g9918,g11279,g10518,g10513,g10440,I16145,g8708,g7055,g5264,g6329,
    g8176,g8005,g7510,g4099,g3281,g11601,g11187,g6746,g6221,g8630,g9622,g11143,
    g10923,g9904,g9886,g9676,g8733,g6624,g11169,g8073,g9841,g9706,g9512,g5882,
    g5592,g8796,g8645,g11168,g4269,g5611,g8069,g9695,g10304,g8469,g8305,g4712,
    g6576,g5762,g10622,g11015,g5217,g5674,g9359,g9173,g9223,g8960,g11556,g9858,
    g5541,g4534,g5897,g6699,g6177,g6855,g3804,g3098,g5680,g9642,g5744,g8399,
    g9447,g9030,g11178,g8510,g8414,g6319,g11186,g3908,g2951,g6352,g9595,g9205,
    g4831,g4109,g5492,g8934,g10312,g6186,g9612,g9417,g9935,g9914,g8701,g10745,
    g10658,g11216,g9328,g8971,g11587,g6325,g7368,g6083,g6544,g5476,g7743,g4869,
    g5722,g6790,g5813,g8408,g10761,g7734,g8136,g7926,g5569,g9902,g9392,g8623,
    g5500,g2496,g6756,g3010,g5877,g8972,g6622,g11612,g9366,g11230,g4364,g9649,
    g5795,g5737,g4054,g6345,g5823,g11275,g9851,g6763,g5802,I16142,g10511,
    g10509,g10507,g9698,g4725,g9964,g9954,g5523,g8550,g8402,g8845,g8611,g2081,
    g6359,g11586,g11007,g5147,g5104,g5099,g4821,g5919,g5499,g4389,g3529,g6416,
    g3497,g4990,g9619,g9010,I6630,g6047,g9652,g10505,g10469,g9843,g9711,g9519,
    g5273,g11465,g4348,g11237,g9834,g9731,g6654,g5444,g3714,g11285,g9598,g8097,
    g8726,g6880,g4816,g3287,g10759,g9938,g9917,g10758,g10652,g9909,g9891,g7127,
    g6663,g11165,g6328,g8401,g11006,g5125,g4865,g4715,g4604,g2325,g5513,g11222,
    g6554,g7732,g9586,g5178,g4401,g4104,g4584,g7472,g11253,g9860,g8703,g11600,
    g9645,g11236,g4162,g3106,g6090,g9691,g11316,g11175,g8068,g9607,g9962,g9952,
    g6348,g9659,g9358,I6316,I6317,g4486,g9587,g8995,g5632,g8965,g4881,g11209,
    g8848,g8715,g4070,g3263,g6463,g8699,g7820,g11021,g5917,g6619,g6318,g6872,
    g11201,g10514,g10489,g4006,g9853,g11274,g8119,g9420,g5233,g7092,g6549,
    g11464,g4487,g2939,g7060,g6739,g5725,g11615,g2544,g11252,g5532,g11153,
    g3771,g9905,g9872,g9680,g7739,g6321,g8386,g8975,g2306,g6625,g7937,g8303,
    g8170,g5706,g2756,g8821,g8643,g10946,g5225,g4169,g5029,g11164,g4007,g4059,
    g4868,g5675,g4718,g10682,g6687,g7704,g4261,g3422,g5745,g8387,g7954,g11283,
    g8461,g8298,g10760,g11480,g6626,g8756,g6341,g10506,g9648,g7453,g5995,g6645,
    g5707,g7548,g11091,g11174,g8403,g8841,g8605,g6879,g8763,g4502,g9839,g9702,
    g9742,g6358,g5841,g5575,g8107,g10240,g11192,g9618,g5539,g8416,g9693,g11553,
    g7557,g5268,g9107,g10633,g7894,g8654,g9621,g6794,g5819,g4883,g3412,g7661,
    g2800,g3389,g3268,g9908,g3429,g6628,g5470,g7526,g2204,g5025,g6204,g4921,
    g4048,g8935,g2525,g9593,g4827,g10701,g10777,g10733,g8130,g9965,g9955,g3684,
    g11213,g5006,g9933,g9912,g8554,g8407,g9641,g6323,g10766,g10646,g6666,g4994,
    g5103,g11592,g3717,g6875,g9658,g6530,g6207,g8199,g7265,g9835,g9735,g6655,
    g3875,g7970,g7384,g5491,g8949,g11152,g9611,g6410,g2804,g10451,g4397,g7224,
    g5398,g5602,g6884,g8698,g8964,g11413,g4950,g5535,g7277,g6772,g8463,g8301,
    g2511,g10728,g6618,g6235,g6355,g4723,g3626,g8720,g6693,g11020,g11583,g8118,
    g8167,g7892,g8652,g5721,g10367,g10362,g9901,g6792,g11282,g7945,g11302,
    g11105,g3634,g8598,g8471,g7140,g9600,g9864,g11613,g5188,g7435,g7876,g4058,
    g6776,g5809,g10301,g4505,g9623,g10739,g11027,g10738,g8687,g8558,g6360,
    g9871,g5108,g11248,g4992,g11552,g9651,g11204,g7824,g5115,g8710,g7102,g9384,
    g2561,g9838,g9700,g9754,g3718,g10661,g10594,g11321,g8879,g7621,g8962,
    g10715,g2272,g8659,g9643,g8957,g5538,g4000,g4126,g4400,g4088,I5886,I5887,
    g6238,g10727,g8174,g5067,g5418,g10297,g6353,g11026,g11212,g6744,g4828,
    g10671,g4383,g2517,g5256,g4297,g4220,g8380,g8252,g7071,g9613,g8933,g5181,
    g7948,g11149,g9862,g11387,g7955,g4161,g11148,g2321,g9712,g8931,g11097,
    g3819,g11104,g2963,g6092,g4999,g7409,g4976,g6858,g4103,I6309,g6580,g5944,
    g5631,g9414,g9660,g9946,g9926,I6331,g9903,g9885,g9673,g10625,g6623,g11228,
    g11011,g6889,g7523,g7822,g8123,g11582,g4316,g3400,g10969,g3625,g5041,g9335,
    g9831,g9727,g9422,g8648,g4588,g8511,g8875,g5168,g7895,g7503,g8655,g3396,
    g4914,g9947,g9927,g5772,g5531,g5036,g10503,g8010,g7738,g8410,g6231,g5608,
    g10581,g10450,g10364,g2132,g2379,g4820,g9653,g10818,g8172,g10429,g5074,
    g9869,g10741,g10635,g8693,g5480,g4581,g3766,g2981,g8555,g8409,g9364,g8994,
    g11299,g6592,g7958,g4995,g4079,g2264,g2160,g3257,I6310,g5000,g3301,I5084,
    g9412,g9389,g10706,g10567,g10366,g10447,g10446,g10533,g5220,g10624,g10300,
    g5023,g4432,g4053,g7596,g5588,g6074,g9963,g9953,g3772,g3089,g5051,g8724,
    g4157,g9707,g8878,g10763,g10639,g6777,g8109,g7898,g7511,g11271,g11461,
    g5732,g11145,g11031,g9865,g9715,g9604,g8799,g8647,g11198,g6873,g6632,g6095,
    g9833,g9729,g6102,g7819,g11280,g7088,g9584,g9896,g8209,g6752,g11161,g8947,
    g5681,g7951,g9419,g5533,g8936,g10670,g11087,g4949,g6364,g5851,g7825,g10667,
    g7136,g6532,g9385,g9897,g9425,g3383,g5601,g7943,g11171,I6631,g7230,g6064,
    g4952,g8736,g6787,g8968,g10306,g11459,g11458,g5739,g7496,g4986,g11010,
    g5187,g3999,g8175,g8722,g5590,g7891,g7471,g8651,g5479,g11599,g6684,g6745,
    g6639,g3696,g4503,g6791,g8180,g4224,g5501,g8838,g8602,g10666,g11158,g9602,
    g5704,g4617,g3879,g9868,g11295,g11144,g9718,g3434,g4987,g6098,g9582,g3533,
    g8104,g9415,g8499,g8377,g9664,g2534,g8754,g9413,g6162,g3584,g4991,g6362,
    g5846,g10685,g11023,g7598,g11224,g11571,g4959,g5626,g9940,g9920,g4876,
    g6730,g9689,g10762,g6070,g9428,g9430,g8927,g7068,g8014,g7740,g11278,g5782,
    g9910,g4236,g11559,g9609,g11558,g6087,g4877,g10751,g10772,g10655,g8135,
    g11544,g5084,g8382,g10230,g7241,g3942,g10638,g4064,g9365,g9861,g9738,g9579,
    g8749,g11255,g11189,g10510,g2917,g11188,g9846,g7818,g11460,g11030,g11093,
    g7893,g7478,g8653,g10442,g6535,g8102,I5085,g3912,g7186,g4489,g9662,g9418,
    g11218,g10746,g10643,g7125,g7821,g6246,g8963,g7533,g10237,g7939,g8786,
    g8638,g10684,g11455,g8364,g2990,g9847,g7584,g5617,g5981,g5789,g4009,g11277,
    g6940,g6472,g7061,g6760,g11595,g5771,g8553,g8405,g4836,g5547,g4967,g6671,
    g7200,g7046,g4229,g8389,g6430,g8706,g4993,g6247,g11170,g7145,g5738,g3998,
    g6741,g11167,g11194,g11589,g4431,g7536,g9585,g2957,g11588,g5690,g6883,
    g4837,g8791,g8641,g6217,g11022,g5915,g4168,g8759,g5110,g11254,g7567,g4392,
    g3273,g9856,g9411,g5002,g11101,g11177,g11560,g8098,g3970,g4941,g6662,g7935,
    g6067,g9863,g9740,g6994,g6758,g4252,g11166,g7130,g11009,g5179,g7542,g11008,
    g5171,g3516,g7573,g3987,g11555,g9857,g9734,g9569,g8728,g8730,g8185,g8385,
    g7902,g4073,g8070,g5731,g11238,g8470,g8308,g5489,g3991,g7823,g4069,g11176,
    g11092,g11154,g9608,g11637,g2091,g8406,g5254,g8612,g9588,g8801,g8742,g7063,
    g10303,g5009,g9665,g8748,g11215,g10750,g5769,g3818,g8755,g6673,g7720,g4609,
    g7547,g7971,g11288,g7599,g6058,g6743,g4106,g6890,g7549,g7269,g8169,g11304,
    g9944,g9924,g7592,g8718,g8616,g9316,g7625,g8793,g8644,g2940,g11624,g10949,
    g2947,g4870,g3563,g10948,g2223,g8246,g7846,g5788,g4008,g9596,g5249,g11585,
    g4972,g11554,g7096,g10673,g4806,g2493,g9936,g9915,g2910,g9317,g10933,
    g10853,g8388,g8177,g7141,g10508,g4230,g10634,g9601,g9192,g6326,g7710,g8028,
    g7375,g5640,g5031,g4550,g7879,g7962,g9597,g5005,g6423,g8108,g5911,g3322,
    g9937,g9916,g9840,g9704,g9747,g10723,g8217,g11013,g5209,g9390,g11214,g6327,
    g5796,g5473,g6346,g5038,g6633,g11005,g5119,g8365,g7558,g4481,g4097,g7588,
    g4497,g9942,g9922,g6696,g10731,g5118,g10665,g8827,g8552,g5540,g4960,g8846,
    g8615,g5983,g6240,g7931,g11100,g11235,g5199,g6316,g7515,g5781,g8018,g7742,
    g2950,g5510,g6347,g9357,g11407,g10743,g5259,g5694,g10769,g11584,g4932,
    g10768,g10649,g4068,g6317,g5215,g4276,g4866,g6775,g10662,g8101,g5825,g3204,
    g5318,g7884,g7457,g3974,g9949,g9929,g10778,g7524,g6079,g7235,g9603,g9850,
    g9726,g9560,g7988,g5228,g5587,g5934,g8168,g9583,g10672,g8627,g8309,g10449,
    g10420,g11273,g8734,g5913,g4572,g6363,g11463,g8074,g8474,g8383,g11234,
    g4483,g11491,g5097,g5726,g5497,g7933,g9617,g9906,g9873,g9683,g11012,g5196,
    g7050,g10971,g10849,g8400,g4345,g9945,g9925,g7271,g5028,g9709,g4223,g10716,
    g10497,g11247,g6661,g11173,g6075,g8023,g7367,g9907,g9888,g9686,g10582,
    g5746,g9959,g9950,g7674,g9690,g5703,g4522,g4115,g7075,g10627,g4047,g2944,
    g6646,g7132,g11029,g7572,g8127,g7209,g11028,g10742,g8880,g10681,g9663,
    g5349,g8732,g3807,g8753,g5848,g3860,g8508,g8411,g8072,g5699,g11240,g6616,
    g6105,g10690,g7582,g9590,g4128,g6404,g6647,g10504,g9657,g4542,g5524,g9899,
    g7736,g10626,g6320,g7623,g10299,g7889,g10298,g8413,g3979,g5211,g4512,g7722,
    g9844,g9714,g9522,g4823,g5993,g5026,g8705,g10737,g10232,g6771,g5170,g8117,
    g9966,g9956,g5280,g7139,g11099,g6892,g9705,g10512,g11098,g8628,g5544,
    g11272,g5483,g9948,g9928,g4063,g11462,g6738,g7593,g11032,g10445,g8882,
    g10316,g5756,g4720,g9409,g8929,g6876,g4989,g9836,g9737,g6061,g8268,g6465,
    g5003,g9967,g9957,g5145,g4834,g4971,g10753,g5695,g7613,g10736,g11220,g7444,
    g4670,g4253,g8163,g7960,g10764,g5757,g10365,g8032,g7385,g11591,g2988,g7583,
    g11147,g5522,g9837,g9697,g9751,g9620,g11151,g11172,g7885,g5595,g5537,g9842,
    g9708,g9516,g4141,g4341,g7679,g7378,g5612,g3939,g7135,g10970,g11025,g9854,
    g9730,g9566,g7182,g9941,g9921,g6194,g4962,g4358,g8683,g4803,g8549,g5224,
    g8778,g11281,g8735,g11146,g3904,g2948,g8075,g9829,g9723,g7184,g11246,g6350,
    g5837,g5902,g2555,g6438,g5512,g5090,g7719,g3695,g7587,g9610,g3536,g8881,
    g4559,g10561,g10549,g5698,g11226,g10295,g5260,g10680,g11551,g11538,g9849,
    g5279,g8404,g5720,g8764,g11318,g11297,g9898,g9510,g7963,g9759,g9803,g6124,
    I14585,I5600,g9489,g3107,g2167,g9362,I14866,g4997,g10291,g9669,g6122,g9509,
    g5227,I15054,g5555,g10376,g8249,I15210,g9882,I5805,g2102,g2099,g2096,g2088,
    I15039,g8259,g10805,I15214,I15215,g8322,g9750,g8248,g8154,I6351,g2405,
    g2389,g2380,g2372,I16427,I14776,g4052,g2862,g2515,I14858,I15209,g2528,
    g2522,g9515,g3118,g2180,I5571,g2514,I5599,g9528,I5629,g2315,I5363,g8159,
    g10521,I16148,I16149,g8417,I14855,I15205,g9878,I15051,g9615,g8823,g8148,
    g2863,g2516,g9511,g9654,I15224,I15225,g8253,g9416,I15171,I15172,g9410,
    I15204,I14596,g9655,g10472,g10470,g10468,g10467,g10386,g10384,g10476,
    g10474,g8158,g9656,g9746,I5357,g9758,I5626,I15057,I15219,I15220,g9616,
    I14862,g2521,I14751,g9591,g9757,g9815,I14835,I16161,g10479,g10478,g10477,
    g10475,g2353,g9776,I5804,I15199,g8153,g9881,g9426,g9423,g8262,g2499,I5570,
    I14607,g9388,g10807,I16160,g10394,g10392,g10482,g10481,I15042,g9589,g9667,
    I14827,g9779,g9391,g2309,I5358,I15177,g9876,g9421,g5186,I6350,g8162,I14779,
    g2305,I5351,I5352,I15176,g9879,g10562,g9606,I14822,I15200,g9880,I14582,
    g8247,I5576,g4476,g2538,I5649,g9605,g9781,g9363,I14831,g8263,g9361,g5780,
    I15048,g9647,g9817,I14602,I15033,g2445,g2437,g2433,g2419,I5366,g9506,g8161,
    g2316,g4675,g9387,I15045,g9808,g2501,g9877,g10529,g9874,g8157,g6899,g9646,
    g2111,g2109,g2106,g2104,I5612,I5613,I5593,I5591,g8970,g8839,I10519,I11279,
    I11278,g3978,I5264,I5263,I8640,g4278,I6761,g2943,I6760,I17400,g11418,
    g11416,I5450,I5449,I16060,g10372,I16058,I6746,g2938,I11975,I11973,I12136,
    I11937,I11935,g2959,I6167,I6168,I5878,g2120,g2115,I5619,I5620,g5552,I6468,
    I6467,I8796,g4672,I8795,I15891,I15892,I5611,g8738,I6716,I6714,I7685,g3460,
    I7683,I12108,I12106,I6747,g2236,I5230,I5231,I12075,I12076,I15870,g10358,
    I16067,I16065,I7562,I13531,I13529,I8797,I17584,I11936,I15257,I15256,I13505,
    I13506,g8824,g8502,g8501,I6186,g11496,I17504,I17505,I16001,I15999,I6125,
    g2215,I6124,I11909,I11907,I12040,I12038,I13909,I13907,I6771,I6772,I11908,
    I16008,I16009,I13908,I7034,I7035,I8650,I9947,I9948,I16066,g10428,I6144,
    I6145,I11242,I11241,I15993,I15994,I6187,g6027,I5500,I11974,I12062,I12060,
    I8771,I8772,I5184,I13293,I6200,I6199,I13265,I5024,I5023,I7863,I13991,
    I13992,I13660,I13661,I6143,I13990,I11510,I11508,g5034,I5229,I12047,I12045,
    I10771,I10769,I16045,I16046,I12061,I5104,I13530,I6447,I4956,I4954,I8481,
    g3530,I8479,I8739,I8740,I6880,I6879,I15431,I15430,I12020,I12019,I16331,
    I16332,I16469,I16467,I5014,I5013,I13523,I13521,I16039,I16037,I16468,I12046,
    I16038,g10427,I8676,g4374,I12113,I8761,g4616,g10422,I15992,I5036,I5034,
    I14263,g8843,I13249,I13250,I5135,I5485,I5486,I7033,I15443,I15441,I6166,
    I8624,g4267,I16015,g10425,I8677,I8576,g4234,I8575,I14613,g9204,I14612,
    I8716,g4601,I8715,I6715,I13514,I13515,I12003,I12002,g2177,I5127,I5128,
    I8577,I17395,g11414,I17393,I11280,I5265,I6989,I6988,I13274,I13272,I10507,
    I5164,I14443,I14444,I9559,I9557,I5592,I13077,I13078,I8717,I5296,I5295,
    I8625,I8626,I4911,I4912,I16000,g10423,I5371,I5185,I5186,I5675,I8544,g4218,
    I8543,I10520,I10521,I5297,I13537,I13283,g4749,I11982,I11980,I8514,g4873,
    I8513,I13091,I13089,I6126,I15908,g10302,I15906,I8763,g8825,g8506,I16007,
    g10424,I5865,g2107,g2105,I5604,I5517,I5518,I6111,I6109,I4929,I4930,I13522,
    I10770,I5539,I5538,I17394,g11415,I13553,I13552,I8642,I17296,I17297,I14278,
    I14279,I4910,I6794,I6792,I5484,I15442,I10931,I10932,I8779,I8780,g2354,
    I15615,g10043,g10153,I17281,I5470,I5468,I11509,I5025,I14272,I14270,I6208,
    I6209,I17290,I17288,I7563,I7564,I5006,I5005,I12128,I12126,I5105,I6323,
    I6322,I12093,I12094,I6666,g2776,I6664,g3623,I6762,I5373,I8529,I8527,I5283,
    I5282,I7224,I7223,I5007,I5459,I17295,I5015,I14264,I14265,I16073,I16072,
    g3205,I8652,I9558,I5203,I5202,I6806,I6807,I6469,I12145,I12143,I12127,
    I13302,I13300,I5502,I9574,I6448,I6449,I8670,I8669,I15453,I15451,I7876,
    I7875,I14203,I14202,I15607,g10149,g10144,I5324,I5325,I8738,g10434,g5859,
    I8606,I8604,I12087,I12085,I13248,I4979,I4980,I12069,I12067,g8942,I12068,
    I17503,I7877,I5165,I6289,I6287,I6777,I8562,I8563,I15890,I13090,g8006,
    g11474,I17460,I17461,I13513,I4986,I4987,I5204,I13504,I6207,I12086,I8545,
    I8180,I8178,I8591,I8589,I10930,I17402,I13294,I13295,I12144,g8757,g2961,
    I14211,I14209,I8515,I5316,I5317,I9946,I8750,g4613,I5605,I14204,I16051,
    g10371,g10373,g10360,g6037,I13858,I13859,I15872,I8528,g4879,I13901,I13902,
    g8542,I6838,I6836,I17307,I17305,g4538,I15452,I13857,I13765,I8671,g10370,
    I16044,g10363,g5360,I5106,I8804,g4677,I8803,I16016,I16017,I17487,I17485,
    I4995,I12092,I8678,I5126,I5372,I17306,I11995,I7225,I11261,g8545,I6110,
    I4942,I4941,I15899,I15900,g5527,g10443,g5350,I16081,g10374,I16079,I8641,
    I6178,I6176,I12074,I5451,I7322,I7323,I6288,I8179,I6805,I17486,I4928,g10286,
    I16330,I9575,I13887,I13886,I8787,I8788,I5315,g10285,I13869,I13867,I13868,
    I13259,I13258,g3261,I16074,I5136,I5137,I5460,I5461,I8605,I6770,g11449,
    I17401,g11448,I15717,g10231,I15716,I14210,I17569,I17567,I13878,I13876,
    I5606,I14442,I11996,I11997,I14277,I17568,I7321,I6990,g8847,I9006,I4985,
    I8651,I13545,I13544,I13894,I13895,I6138,I6136,I13076,g2205,I13260,I5501,
    I17586,I13900,I6201,I14217,g8826,I14216,I9007,I13561,I13559,g10229,I17493,
    I17492,I12215,I12214,I11262,I11263,I6225,I6226,I13309,I13307,I5676,I5677,
    I6826,I6827,I13308,g8190,g2792,I5879,I5880,g3061,I17585,I6881,I12138,I8729,
    g4605,I8728,I15871,I5866,I5867,I6793,I6487,I16080,I13893,I12115,I6748,
    I6224,I8805,I15880,I15878,I16031,I16030,I14271,I13267,I15616,I15617,I4966,
    I4964,I8752,I15432,g10438,g6032,g3011,I8480,I16087,I16086,g3734,I14218,
    I4955,I8786,g4639,g10480,I11915,I11914,I8770,g4619,I5516,g8541,I6188,I5892,
    I5891,I13766,I13767,I15258,I13266,I6825,I17283,g5277,I5035,g10375,I15879,
    g10359,I12114,I12107,g2500,g10430,g5999,I13285,I13877,g2795,I5893,I13560,
    g4259,I5166,I14614,I4965,I4943,I16023,g10426,I16059,g8737,I9576,I16052,
    I16053,I12004,g5573,I6837,I8730,I4978,I6177,I17051,I7864,I7865,I6665,
    I12216,I13554,g10368,I13284,I6137,I5529,I5530,I17282,I5618,I8664,I8662,
    I11916,g7717,I4972,I4971,I13273,I10509,I10508,I6778,I6779,I5469,g4251,
    I13546,I4996,I4997,I13539,I16032,I5323,I13538,I5540,I8778,g4286,I17052,
    I17053,g10287,I15898,g7978,g4227,I8561,I8762,I8751,I15907,I4973,I16024,
    I16025,g4455,I5342,I5341,I12137,g10483,I16088,I17289,g4630,I15609,I15608,
    g10436,g6023,I17459,I13301,I11981,I8663,I15718,I5284,g4607,g8840,g10441,
    g5345,g10432,g5938,I12021,I6489,I5528,I13659,I5343,I12039,I9008,I6488,
    I13888,I17494,I7684,g3221,I6324,I8590,I11243,g10324,g10239,g4974,g10322;

  FD1 DFF_0(CK,g1289,g5660);
  FD1 DFF_1(CK,g1882,g9349);
  FD1 DFF_2(CK,g312,g5644);
  FD1 DFF_3(CK,g452,g11257);
  FD1 DFF_4(CK,g123,g8272);
  FD1 DFF_5(CK,g207,g7315);
  FD1 DFF_6(CK,g713,g9345);
  FD1 DFF_7(CK,g1153,g6304);
  FD1 DFF_8(CK,g1209,g10873);
  FD1 DFF_9(CK,g1744,g5663);
  FD1 DFF_10(CK,g1558,g7349);
  FD1 DFF_11(CK,g695,g9343);
  FD1 DFF_12(CK,g461,g11467);
  FD1 DFF_13(CK,g940,g8572);
  FD1 DFF_14(CK,g976,g11471);
  FD1 DFF_15(CK,g709,g8432);
  FD1 DFF_16(CK,g1092,g6810);
  FD1 DFF_17(CK,g1574,g7354);
  FD1 DFF_18(CK,g1864,g7816);
  FD1 DFF_19(CK,g369,g11439);
  FD1 DFF_20(CK,g1580,g7356);
  FD1 DFF_21(CK,g1736,g6846);
  FD1 DFF_22(CK,g39,g10774);
  FD1 DFF_23(CK,g1651,g11182);
  FD1 DFF_24(CK,g1424,g7330);
  FD1 DFF_25(CK,g1737,g1736);
  FD1 DFF_26(CK,g1672,g11037);
  FD1 DFF_27(CK,g1077,g6805);
  FD1 DFF_28(CK,g1231,g8279);
  FD1 DFF_29(CK,g4,g8079);
  FD1 DFF_30(CK,g774,g7785);
  FD1 DFF_31(CK,g1104,g6815);
  FD1 DFF_32(CK,g1304,g7290);
  FD1 DFF_33(CK,g243,g7325);
  FD1 DFF_34(CK,g1499,g8447);
  FD1 DFF_35(CK,g1044,g7789);
  FD1 DFF_36(CK,g1444,g8987);
  FD1 DFF_37(CK,g757,g11179);
  FD1 DFF_38(CK,g786,g8436);
  FD1 DFF_39(CK,g1543,g7344);
  FD1 DFF_40(CK,g552,g11045);
  FD1 DFF_41(CK,g315,g5645);
  FD1 DFF_42(CK,g1534,g7341);
  FD1 DFF_43(CK,g622,g9338);
  FD1 DFF_44(CK,g1927,g9354);
  FD1 DFF_45(CK,g1660,g11033);
  FD1 DFF_46(CK,g278,g7765);
  FD1 DFF_47(CK,g1436,g8989);
  FD1 DFF_48(CK,g718,g8433);
  FD1 DFF_49(CK,g76,g7775);
  FD1 DFF_50(CK,g554,g11047);
  FD1 DFF_51(CK,g496,g11333);
  FD1 DFF_52(CK,g981,g11472);
  FD1 DFF_53(CK,g878,g4896);
  FD1 DFF_54(CK,g590,g5653);
  FD1 DFF_55(CK,g829,g4182);
  FD1 DFF_56(CK,g1095,g6811);
  FD1 DFF_57(CK,g704,g9344);
  FD1 DFF_58(CK,g1265,g7302);
  FD1 DFF_59(CK,g1786,g7814);
  FD1 DFF_60(CK,g682,g8429);
  FD1 DFF_61(CK,g1296,g7292);
  FD1 DFF_62(CK,g587,g6295);
  FD1 DFF_63(CK,g52,g7777);
  FD1 DFF_64(CK,g646,g8065);
  FD1 DFF_65(CK,g327,g5649);
  FD1 DFF_66(CK,g1389,g6836);
  FD1 DFF_67(CK,g1371,g7311);
  FD1 DFF_68(CK,g1956,g1955);
  FD1 DFF_69(CK,g1675,g11038);
  FD1 DFF_70(CK,g354,g11508);
  FD1 DFF_71(CK,g113,g7285);
  FD1 DFF_72(CK,g639,g8063);
  FD1 DFF_73(CK,g1684,g11041);
  FD1 DFF_74(CK,g1639,g8448);
  FD1 DFF_75(CK,g1791,g8080);
  FD1 DFF_76(CK,g248,g7323);
  FD1 DFF_77(CK,g1707,g4907);
  FD1 DFF_78(CK,g1759,g5668);
  FD1 DFF_79(CK,g351,g11507);
  FD1 DFF_80(CK,g1957,g1956);
  FD1 DFF_81(CK,g1604,g7364);
  FD1 DFF_82(CK,g1098,g6812);
  FD1 DFF_83(CK,g932,g8570);
  FD1 DFF_84(CK,g126,g5642);
  FD1 DFF_85(CK,g1896,g8282);
  FD1 DFF_86(CK,g736,g8435);
  FD1 DFF_87(CK,g1019,g7807);
  FD1 DFF_88(CK,g1362,g7305);
  FD1 DFF_89(CK,g745,g2639);
  FD1 DFF_90(CK,g1419,g7332);
  FD1 DFF_91(CK,g58,g7779);
  FD1 DFF_92(CK,g32,g11397);
  FD1 DFF_93(CK,g876,g878);
  FD1 DFF_94(CK,g1086,g6808);
  FD1 DFF_95(CK,g1486,g8444);
  FD1 DFF_96(CK,g1730,g10881);
  FD1 DFF_97(CK,g1504,g7328);
  FD1 DFF_98(CK,g1470,g8440);
  FD1 DFF_99(CK,g822,g8437);
  FD1 DFF_100(CK,g583,g6291);
  FD1 DFF_101(CK,g1678,g11039);
  FD1 DFF_102(CK,g174,g8423);
  FD1 DFF_103(CK,g1766,g7810);
  FD1 DFF_104(CK,g1801,g8450);
  FD1 DFF_105(CK,g186,g7317);
  FD1 DFF_106(CK,g959,g11403);
  FD1 DFF_107(CK,g1169,g6314);
  FD1 DFF_108(CK,g1007,g7806);
  FD1 DFF_109(CK,g1407,g8993);
  FD1 DFF_110(CK,g1059,g7794);
  FD1 DFF_111(CK,g1868,g7817);
  FD1 DFF_112(CK,g758,g6797);
  FD1 DFF_113(CK,g1718,g6337);
  FD1 DFF_114(CK,g396,g11265);
  FD1 DFF_115(CK,g1015,g7808);
  FD1 DFF_116(CK,g38,g10872);
  FD1 DFF_117(CK,g632,g5655);
  FD1 DFF_118(CK,g1415,g7335);
  FD1 DFF_119(CK,g1227,g8278);
  FD1 DFF_120(CK,g1721,g10878);
  FD1 DFF_121(CK,g882,g883);
  FD1 DFF_122(CK,g16,g4906);
  FD1 DFF_123(CK,g284,g7767);
  FD1 DFF_124(CK,g426,g11256);
  FD1 DFF_125(CK,g219,g7310);
  FD1 DFF_126(CK,g1216,g1360);
  FD1 DFF_127(CK,g806,g7289);
  FD1 DFF_128(CK,g1428,g8992);
  FD1 DFF_129(CK,g579,g6287);
  FD1 DFF_130(CK,g1564,g7351);
  FD1 DFF_131(CK,g1741,g5662);
  FD1 DFF_132(CK,g225,g7309);
  FD1 DFF_133(CK,g281,g7766);
  FD1 DFF_134(CK,g1308,g11627);
  FD1 DFF_135(CK,g611,g9930);
  FD1 DFF_136(CK,g631,g5654);
  FD1 DFF_137(CK,g1217,g9823);
  FD1 DFF_138(CK,g1589,g7359);
  FD1 DFF_139(CK,g1466,g8439);
  FD1 DFF_140(CK,g1571,g7353);
  FD1 DFF_141(CK,g1861,g7815);
  FD1 DFF_142(CK,g1365,g7307);
  FD1 DFF_143(CK,g1448,g11594);
  FD1 DFF_144(CK,g1711,g6335);
  FD1 DFF_145(CK,g1133,g6309);
  FD1 DFF_146(CK,g1333,g11635);
  FD1 DFF_147(CK,g153,g8426);
  FD1 DFF_148(CK,g962,g11404);
  FD1 DFF_149(CK,g766,g6799);
  FD1 DFF_150(CK,g588,g6296);
  FD1 DFF_151(CK,g486,g11331);
  FD1 DFF_152(CK,g471,g11469);
  FD1 DFF_153(CK,g1397,g7322);
  FD1 DFF_154(CK,g580,g6288);
  FD1 DFF_155(CK,g1950,g8288);
  FD1 DFF_156(CK,g756,g755);
  FD1 DFF_157(CK,g635,g5656);
  FD1 DFF_158(CK,g1101,g6814);
  FD1 DFF_159(CK,g549,g11044);
  FD1 DFF_160(CK,g1041,g7788);
  FD1 DFF_161(CK,g105,g11180);
  FD1 DFF_162(CK,g1669,g11036);
  FD1 DFF_163(CK,g1368,g7308);
  FD1 DFF_164(CK,g1531,g7340);
  FD1 DFF_165(CK,g1458,g7327);
  FD1 DFF_166(CK,g572,g10877);
  FD1 DFF_167(CK,g1011,g7805);
  FD1 DFF_168(CK,g33,g10867);
  FD1 DFF_169(CK,g1411,g7331);
  FD1 DFF_170(CK,g1074,g6813);
  FD1 DFF_171(CK,g444,g11259);
  FD1 DFF_172(CK,g1474,g8441);
  FD1 DFF_173(CK,g1080,g6806);
  FD1 DFF_174(CK,g1713,g6336);
  FD1 DFF_175(CK,g333,g5651);
  FD1 DFF_176(CK,g269,g7762);
  FD1 DFF_177(CK,g401,g11266);
  FD1 DFF_178(CK,g1857,g11409);
  FD1 DFF_179(CK,g9,g7336);
  FD1 DFF_180(CK,g664,g8782);
  FD1 DFF_181(CK,g965,g11405);
  FD1 DFF_182(CK,g1400,g7324);
  FD1 DFF_183(CK,g309,g5652);
  FD1 DFF_184(CK,g814,g8077);
  FD1 DFF_185(CK,g231,g7319);
  FD1 DFF_186(CK,g557,g11048);
  FD1 DFF_187(CK,g586,g6294);
  FD1 DFF_188(CK,g869,g875);
  FD1 DFF_189(CK,g1383,g7316);
  FD1 DFF_190(CK,g158,g8425);
  FD1 DFF_191(CK,g627,g5657);
  FD1 DFF_192(CK,g1023,g7799);
  FD1 DFF_193(CK,g259,g7755);
  FD1 DFF_194(CK,g1361,g1206);
  FD1 DFF_195(CK,g1327,g11633);
  FD1 DFF_196(CK,g654,g8067);
  FD1 DFF_197(CK,g293,g7770);
  FD1 DFF_198(CK,g1346,g11656);
  FD1 DFF_199(CK,g1633,g8873);
  FD1 DFF_200(CK,g1753,g5666);
  FD1 DFF_201(CK,g1508,g7329);
  FD1 DFF_202(CK,g1240,g7297);
  FD1 DFF_203(CK,g538,g11326);
  FD1 DFF_204(CK,g416,g11269);
  FD1 DFF_205(CK,g542,g11325);
  FD1 DFF_206(CK,g1681,g11040);
  FD1 DFF_207(CK,g374,g11440);
  FD1 DFF_208(CK,g563,g11050);
  FD1 DFF_209(CK,g1914,g8284);
  FD1 DFF_210(CK,g530,g11328);
  FD1 DFF_211(CK,g575,g11052);
  FD1 DFF_212(CK,g1936,g9355);
  FD1 DFF_213(CK,g55,g7778);
  FD1 DFF_214(CK,g1117,g6299);
  FD1 DFF_215(CK,g1317,g1356);
  FD1 DFF_216(CK,g357,g11509);
  FD1 DFF_217(CK,g386,g11263);
  FD1 DFF_218(CK,g1601,g7363);
  FD1 DFF_219(CK,g553,g11046);
  FD1 DFF_220(CK,g166,g7747);
  FD1 DFF_221(CK,g501,g11334);
  FD1 DFF_222(CK,g262,g7758);
  FD1 DFF_223(CK,g1840,g8694);
  FD1 DFF_224(CK,g70,g7783);
  FD1 DFF_225(CK,g318,g5646);
  FD1 DFF_226(CK,g1356,g6818);
  FD1 DFF_227(CK,g794,g6800);
  FD1 DFF_228(CK,g36,g10870);
  FD1 DFF_229(CK,g302,g7773);
  FD1 DFF_230(CK,g342,g11513);
  FD1 DFF_231(CK,g1250,g7299);
  FD1 DFF_232(CK,g1163,g6301);
  FD1 DFF_233(CK,g1810,g2044);
  FD1 DFF_234(CK,g1032,g7800);
  FD1 DFF_235(CK,g1432,g8990);
  FD1 DFF_236(CK,g1053,g7792);
  FD1 DFF_237(CK,g1453,g7326);
  FD1 DFF_238(CK,g363,g11511);
  FD1 DFF_239(CK,g330,g5650);
  FD1 DFF_240(CK,g1157,g6303);
  FD1 DFF_241(CK,g1357,g6330);
  FD1 DFF_242(CK,g35,g10869);
  FD1 DFF_243(CK,g928,g8569);
  FD1 DFF_244(CK,g261,g7757);
  FD1 DFF_245(CK,g516,g11337);
  FD1 DFF_246(CK,g254,g7759);
  FD1 DFF_247(CK,g778,g8076);
  FD1 DFF_248(CK,g861,g4190);
  FD1 DFF_249(CK,g1627,g8871);
  FD1 DFF_250(CK,g1292,g7293);
  FD1 DFF_251(CK,g290,g7769);
  FD1 DFF_252(CK,g1850,g5671);
  FD1 DFF_253(CK,g770,g7288);
  FD1 DFF_254(CK,g1583,g7357);
  FD1 DFF_255(CK,g466,g11468);
  FD1 DFF_256(CK,g1561,g7350);
  FD1 DFF_257(CK,g1527,g4899);
  FD1 DFF_258(CK,g1546,g7345);
  FD1 DFF_259(CK,g287,g7768);
  FD1 DFF_260(CK,g560,g11049);
  FD1 DFF_261(CK,g617,g8780);
  FD1 DFF_262(CK,g17,g4894);
  FD1 DFF_263(CK,g336,g11653);
  FD1 DFF_264(CK,g456,g11466);
  FD1 DFF_265(CK,g305,g5643);
  FD1 DFF_266(CK,g345,g11642);
  FD1 DFF_267(CK,g8,g2613);
  FD1 DFF_268(CK,g1771,g7811);
  FD1 DFF_269(CK,g865,g8275);
  FD1 DFF_270(CK,g255,g7751);
  FD1 DFF_271(CK,g1945,g9356);
  FD1 DFF_272(CK,g1738,g5661);
  FD1 DFF_273(CK,g1478,g8442);
  FD1 DFF_274(CK,g1035,g7787);
  FD1 DFF_275(CK,g1959,g4217);
  FD1 DFF_276(CK,g1690,g6844);
  FD1 DFF_277(CK,g1482,g8443);
  FD1 DFF_278(CK,g1110,g6817);
  FD1 DFF_279(CK,g296,g7771);
  FD1 DFF_280(CK,g1663,g11034);
  FD1 DFF_281(CK,g700,g8431);
  FD1 DFF_282(CK,g1762,g5669);
  FD1 DFF_283(CK,g360,g11510);
  FD1 DFF_284(CK,g192,g6837);
  FD1 DFF_285(CK,g1657,g10875);
  FD1 DFF_286(CK,g722,g9346);
  FD1 DFF_287(CK,g61,g7780);
  FD1 DFF_288(CK,g566,g11051);
  FD1 DFF_289(CK,g1394,g7809);
  FD1 DFF_290(CK,g1089,g6809);
  FD1 DFF_291(CK,g883,g4897);
  FD1 DFF_292(CK,g1071,g6804);
  FD1 DFF_293(CK,g986,g11473);
  FD1 DFF_294(CK,g971,g11470);
  FD1 DFF_295(CK,g1955,g6338);
  FD1 DFF_296(CK,g143,g7746);
  FD1 DFF_297(CK,g1814,g9825);
  FD1 DFF_298(CK,g1038,g7797);
  FD1 DFF_299(CK,g1212,g1217);
  FD1 DFF_300(CK,g1918,g9353);
  FD1 DFF_301(CK,g782,g8273);
  FD1 DFF_302(CK,g1822,g9826);
  FD1 DFF_303(CK,g237,g7306);
  FD1 DFF_304(CK,g746,g2638);
  FD1 DFF_305(CK,g1062,g7795);
  FD1 DFF_306(CK,g1462,g8438);
  FD1 DFF_307(CK,g178,g7748);
  FD1 DFF_308(CK,g366,g11512);
  FD1 DFF_309(CK,g837,g4184);
  FD1 DFF_310(CK,g599,g9819);
  FD1 DFF_311(CK,g1854,g11408);
  FD1 DFF_312(CK,g944,g11398);
  FD1 DFF_313(CK,g1941,g8287);
  FD1 DFF_314(CK,g170,g8422);
  FD1 DFF_315(CK,g1520,g7334);
  FD1 DFF_316(CK,g686,g9342);
  FD1 DFF_317(CK,g953,g11401);
  FD1 DFF_318(CK,g1958,g6339);
  FD1 DFF_319(CK,g40,g10775);
  FD1 DFF_320(CK,g1765,g3329);
  FD1 DFF_321(CK,g1733,g10882);
  FD1 DFF_322(CK,g1270,g7303);
  FD1 DFF_323(CK,g1610,g6845);
  FD1 DFF_324(CK,g1796,g8280);
  FD1 DFF_325(CK,g1324,g11632);
  FD1 DFF_326(CK,g1540,g7343);
  FD1 DFF_327(CK,g1377,g7312);
  FD1 DFF_328(CK,g1206,g4898);
  FD1 DFF_329(CK,g491,g11332);
  FD1 DFF_330(CK,g1849,g5670);
  FD1 DFF_331(CK,g213,g7313);
  FD1 DFF_332(CK,g1781,g7813);
  FD1 DFF_333(CK,g1900,g9351);
  FD1 DFF_334(CK,g1245,g7298);
  FD1 DFF_335(CK,g108,g11593);
  FD1 DFF_336(CK,g630,g7287);
  FD1 DFF_337(CK,g148,g8427);
  FD1 DFF_338(CK,g833,g4183);
  FD1 DFF_339(CK,g1923,g8285);
  FD1 DFF_340(CK,g936,g8571);
  FD1 DFF_341(CK,g1215,g6315);
  FD1 DFF_342(CK,g1314,g11629);
  FD1 DFF_343(CK,g849,g4187);
  FD1 DFF_344(CK,g1336,g11654);
  FD1 DFF_345(CK,g272,g7763);
  FD1 DFF_346(CK,g1806,g8573);
  FD1 DFF_347(CK,g826,g8568);
  FD1 DFF_348(CK,g1065,g7796);
  FD1 DFF_349(CK,g1887,g8281);
  FD1 DFF_350(CK,g37,g10871);
  FD1 DFF_351(CK,g968,g11406);
  FD1 DFF_352(CK,g1845,g5673);
  FD1 DFF_353(CK,g1137,g6310);
  FD1 DFF_354(CK,g1891,g9350);
  FD1 DFF_355(CK,g1255,g7300);
  FD1 DFF_356(CK,g257,g7753);
  FD1 DFF_357(CK,g874,g9821);
  FD1 DFF_358(CK,g591,g9818);
  FD1 DFF_359(CK,g731,g9347);
  FD1 DFF_360(CK,g636,g8781);
  FD1 DFF_361(CK,g1218,g8276);
  FD1 DFF_362(CK,g605,g9820);
  FD1 DFF_363(CK,g79,g7776);
  FD1 DFF_364(CK,g182,g7749);
  FD1 DFF_365(CK,g950,g11400);
  FD1 DFF_366(CK,g1129,g6308);
  FD1 DFF_367(CK,g857,g4189);
  FD1 DFF_368(CK,g448,g11258);
  FD1 DFF_369(CK,g1828,g9827);
  FD1 DFF_370(CK,g1727,g10880);
  FD1 DFF_371(CK,g1592,g7360);
  FD1 DFF_372(CK,g1703,g6843);
  FD1 DFF_373(CK,g1932,g8286);
  FD1 DFF_374(CK,g1624,g8870);
  FD1 DFF_375(CK,g26,g4885);
  FD1 DFF_376(CK,g1068,g6803);
  FD1 DFF_377(CK,g578,g6286);
  FD1 DFF_378(CK,g440,g11260);
  FD1 DFF_379(CK,g476,g11338);
  FD1 DFF_380(CK,g119,g7745);
  FD1 DFF_381(CK,g668,g9340);
  FD1 DFF_382(CK,g139,g8418);
  FD1 DFF_383(CK,g1149,g6305);
  FD1 DFF_384(CK,g34,g10868);
  FD1 DFF_385(CK,g1848,g7366);
  FD1 DFF_386(CK,g263,g7760);
  FD1 DFF_387(CK,g818,g8274);
  FD1 DFF_388(CK,g1747,g5664);
  FD1 DFF_389(CK,g802,g6802);
  FD1 DFF_390(CK,g275,g7764);
  FD1 DFF_391(CK,g1524,g7338);
  FD1 DFF_392(CK,g1577,g7355);
  FD1 DFF_393(CK,g810,g7786);
  FD1 DFF_394(CK,g391,g11264);
  FD1 DFF_395(CK,g658,g9339);
  FD1 DFF_396(CK,g1386,g7318);
  FD1 DFF_397(CK,g253,g7750);
  FD1 DFF_398(CK,g875,g9822);
  FD1 DFF_399(CK,g1125,g6307);
  FD1 DFF_400(CK,g201,g7304);
  FD1 DFF_401(CK,g1280,g7295);
  FD1 DFF_402(CK,g1083,g6807);
  FD1 DFF_403(CK,g650,g8066);
  FD1 DFF_404(CK,g1636,g8874);
  FD1 DFF_405(CK,g853,g4188);
  FD1 DFF_406(CK,g421,g11270);
  FD1 DFF_407(CK,g762,g6798);
  FD1 DFF_408(CK,g956,g11402);
  FD1 DFF_409(CK,g378,g11441);
  FD1 DFF_410(CK,g1756,g5667);
  FD1 DFF_411(CK,g589,g6297);
  FD1 DFF_412(CK,g841,g4185);
  FD1 DFF_413(CK,g1027,g7798);
  FD1 DFF_414(CK,g1003,g7803);
  FD1 DFF_415(CK,g1403,g8991);
  FD1 DFF_416(CK,g1145,g6312);
  FD1 DFF_417(CK,g1107,g6816);
  FD1 DFF_418(CK,g1223,g8277);
  FD1 DFF_419(CK,g406,g11267);
  FD1 DFF_420(CK,g1811,g11185);
  FD1 DFF_421(CK,g1642,g11183);
  FD1 DFF_422(CK,g1047,g7790);
  FD1 DFF_423(CK,g1654,g10874);
  FD1 DFF_424(CK,g197,g6835);
  FD1 DFF_425(CK,g1595,g7361);
  FD1 DFF_426(CK,g1537,g7342);
  FD1 DFF_427(CK,g727,g8434);
  FD1 DFF_428(CK,g999,g7804);
  FD1 DFF_429(CK,g798,g6801);
  FD1 DFF_430(CK,g481,g11324);
  FD1 DFF_431(CK,g754,g4895);
  FD1 DFF_432(CK,g1330,g11634);
  FD1 DFF_433(CK,g845,g4186);
  FD1 DFF_434(CK,g790,g8567);
  FD1 DFF_435(CK,g1512,g8449);
  FD1 DFF_436(CK,g114,g113);
  FD1 DFF_437(CK,g1490,g8445);
  FD1 DFF_438(CK,g1166,g6300);
  FD1 DFF_439(CK,g1056,g7793);
  FD1 DFF_440(CK,g348,g11506);
  FD1 DFF_441(CK,g868,g874);
  FD1 DFF_442(CK,g1260,g7301);
  FD1 DFF_443(CK,g260,g7756);
  FD1 DFF_444(CK,g131,g8420);
  FD1 DFF_445(CK,g7,g2731);
  FD1 DFF_446(CK,g258,g7754);
  FD1 DFF_447(CK,g521,g11330);
  FD1 DFF_448(CK,g1318,g11630);
  FD1 DFF_449(CK,g1872,g9348);
  FD1 DFF_450(CK,g677,g9341);
  FD1 DFF_451(CK,g582,g6290);
  FD1 DFF_452(CK,g1393,g7320);
  FD1 DFF_453(CK,g1549,g7346);
  FD1 DFF_454(CK,g947,g11399);
  FD1 DFF_455(CK,g1834,g9895);
  FD1 DFF_456(CK,g1598,g7362);
  FD1 DFF_457(CK,g1121,g6306);
  FD1 DFF_458(CK,g1321,g11631);
  FD1 DFF_459(CK,g506,g11335);
  FD1 DFF_460(CK,g546,g11043);
  FD1 DFF_461(CK,g1909,g9352);
  FD1 DFF_462(CK,g755,g6298);
  FD1 DFF_463(CK,g1552,g7347);
  FD1 DFF_464(CK,g584,g6292);
  FD1 DFF_465(CK,g1687,g11042);
  FD1 DFF_466(CK,g1586,g7358);
  FD1 DFF_467(CK,g324,g5648);
  FD1 DFF_468(CK,g1141,g6311);
  FD1 DFF_469(CK,g1570,g4900);
  FD1 DFF_470(CK,g1341,g11655);
  FD1 DFF_471(CK,g1710,g4901);
  FD1 DFF_472(CK,g1645,g11184);
  FD1 DFF_473(CK,g115,g7321);
  FD1 DFF_474(CK,g135,g8419);
  FD1 DFF_475(CK,g525,g11329);
  FD1 DFF_476(CK,g581,g6289);
  FD1 DFF_477(CK,g1607,g7365);
  FD1 DFF_478(CK,g321,g5647);
  FD1 DFF_479(CK,g67,g7782);
  FD1 DFF_480(CK,g1275,g11443);
  FD1 DFF_481(CK,g1311,g11628);
  FD1 DFF_482(CK,g1615,g8868);
  FD1 DFF_483(CK,g382,g11442);
  FD1 DFF_484(CK,g1374,g6825);
  FD1 DFF_485(CK,g266,g7761);
  FD1 DFF_486(CK,g1284,g7294);
  FD1 DFF_487(CK,g1380,g7314);
  FD1 DFF_488(CK,g673,g8428);
  FD1 DFF_489(CK,g1853,g5672);
  FD1 DFF_490(CK,g162,g8424);
  FD1 DFF_491(CK,g411,g11268);
  FD1 DFF_492(CK,g431,g11262);
  FD1 DFF_493(CK,g1905,g8283);
  FD1 DFF_494(CK,g1515,g7333);
  FD1 DFF_495(CK,g1630,g8872);
  FD1 DFF_496(CK,g49,g7774);
  FD1 DFF_497(CK,g991,g7802);
  FD1 DFF_498(CK,g1300,g7291);
  FD1 DFF_499(CK,g339,g11505);
  FD1 DFF_500(CK,g256,g7752);
  FD1 DFF_501(CK,g1750,g5665);
  FD1 DFF_502(CK,g585,g6293);
  FD1 DFF_503(CK,g1440,g8988);
  FD1 DFF_504(CK,g1666,g11035);
  FD1 DFF_505(CK,g1528,g7339);
  FD1 DFF_506(CK,g1351,g11657);
  FD1 DFF_507(CK,g1648,g11181);
  FD1 DFF_508(CK,g127,g8421);
  FD1 DFF_509(CK,g1618,g11611);
  FD1 DFF_510(CK,g1235,g7296);
  FD1 DFF_511(CK,g299,g7772);
  FD1 DFF_512(CK,g435,g11261);
  FD1 DFF_513(CK,g64,g7781);
  FD1 DFF_514(CK,g1555,g7348);
  FD1 DFF_515(CK,g995,g7801);
  FD1 DFF_516(CK,g1621,g8869);
  FD1 DFF_517(CK,g1113,g6313);
  FD1 DFF_518(CK,g643,g8064);
  FD1 DFF_519(CK,g1494,g8446);
  FD1 DFF_520(CK,g1567,g7352);
  FD1 DFF_521(CK,g691,g8430);
  FD1 DFF_522(CK,g534,g11327);
  FD1 DFF_523(CK,g1776,g7812);
  FD1 DFF_524(CK,g569,g10876);
  FD1 DFF_525(CK,g1160,g6302);
  FD1 DFF_526(CK,g1360,g9824);
  FD1 DFF_527(CK,g1050,g7791);
  FD1 DFF_528(CK,g1,g8078);
  FD1 DFF_529(CK,g511,g11336);
  FD1 DFF_530(CK,g1724,g10879);
  FD1 DFF_531(CK,g12,g7337);
  FD1 DFF_532(CK,g1878,g8695);
  FD1 DFF_533(CK,g73,g7784);
  IV  NOT_0(I8854,g4500);
  IV  NOT_1(g5652,I9117);
  IV  NOT_2(I12913,g7845);
  IV  NOT_3(g11354,I17179);
  IV  NOT_4(g6837,I10891);
  IV  NOT_5(I10941,g6555);
  IV  NOT_6(I6979,g2888);
  IV  NOT_7(g5843,I9458);
  IV  NOT_8(g2771,I5854);
  IV  NOT_9(g3537,g3164);
  IV  NOT_10(g6062,I9699);
  IV  NOT_11(I9984,g5529);
  IV  NOT_12(I14382,g8886);
  IV  NOT_13(g7706,I12335);
  IV  NOT_14(I13618,g8345);
  IV  NOT_15(I15181,g9968);
  IV  NOT_16(g6620,I10573);
  IV  NOT_17(I12436,g7659);
  IV  NOT_18(g5193,g4682);
  IV  NOT_19(g6462,I10394);
  IV  NOT_20(g8925,I14252);
  IV  NOT_21(I14519,g9106);
  IV  NOT_22(g10289,I15691);
  IV  NOT_23(I14176,g8784);
  IV  NOT_24(I14185,g8790);
  IV  NOT_25(g11181,I16944);
  IV  NOT_26(I14675,g9263);
  IV  NOT_27(g2299,g1707);
  IV  NOT_28(I12607,g7633);
  IV  NOT_29(g3272,g2450);
  IV  NOT_30(g2547,g23);
  IV  NOT_31(g9291,g8892);
  IV  NOT_32(I6001,g2548);
  IV  NOT_33(I7048,g2807);
  IV  NOT_34(g10309,I15733);
  IV  NOT_35(g7029,I11180);
  IV  NOT_36(g4440,g4130);
  IV  NOT_37(I9544,g5024);
  IV  NOT_38(g10288,I15688);
  IV  NOT_39(I12274,g7110);
  IV  NOT_40(I9483,g5050);
  IV  NOT_41(g7787,I12526);
  IV  NOT_42(I6676,g2759);
  IV  NOT_43(I8520,g4338);
  IV  NOT_44(g10571,I16236);
  IV  NOT_45(I17692,g11596);
  IV  NOT_46(I17761,g11652);
  IV  NOT_47(I13469,g8147);
  IV  NOT_48(g9344,I14537);
  IV  NOT_49(g7956,g7432);
  IV  NOT_50(g3417,I6624);
  IV  NOT_51(g4323,g4130);
  IV  NOT_52(I11286,g6551);
  IV  NOT_53(I8031,g3540);
  IV  NOT_54(g7675,I12300);
  IV  NOT_55(g8320,I13344);
  IV  NOT_56(I12565,g7388);
  IV  NOT_57(I16644,g10865);
  IV  NOT_58(I11306,g6731);
  IV  NOT_59(g1981,g650);
  IV  NOT_60(I7333,g3729);
  IV  NOT_61(I13039,g8054);
  IV  NOT_62(g3982,g3052);
  IV  NOT_63(g6249,I10006);
  IV  NOT_64(g9259,g8892);
  IV  NOT_65(I15190,g9974);
  IV  NOT_66(g11426,I17331);
  IV  NOT_67(g9819,I14958);
  IV  NOT_68(g8277,I13203);
  IV  NOT_69(I5050,g1216);
  IV  NOT_70(I5641,g546);
  IV  NOT_71(g5121,g4682);
  IV  NOT_72(g1997,g798);
  IV  NOT_73(g3629,g3228);
  IV  NOT_74(g3328,I6501);
  IV  NOT_75(I12641,g7709);
  IV  NOT_76(g5670,I9171);
  IV  NOT_77(g6842,I10898);
  IV  NOT_78(g8617,g8465);
  IV  NOT_79(I15520,g10035);
  IV  NOT_80(I7396,g4102);
  IV  NOT_81(I7803,g3820);
  IV  NOT_82(g3330,I6507);
  IV  NOT_83(g2991,I6233);
  IV  NOT_84(I9461,g4940);
  IV  NOT_85(g2244,I5251);
  IV  NOT_86(g6192,I9923);
  IV  NOT_87(g6298,I10153);
  IV  NOT_88(g6085,I9734);
  IV  NOT_89(I12153,g6874);
  IV  NOT_90(g4351,I7630);
  IV  NOT_91(I11677,g7056);
  IV  NOT_92(g10687,I16356);
  IV  NOT_93(g4530,I7935);
  IV  NOT_94(g8516,I13717);
  IV  NOT_95(g5232,g4640);
  IV  NOT_96(I13975,g8588);
  IV  NOT_97(g2078,g135);
  IV  NOT_98(I8911,g4565);
  IV  NOT_99(g2340,g1918);
  IV  NOT_100(g7684,g7148);
  IV  NOT_101(I12409,g7501);
  IV  NOT_102(g7745,I12400);
  IV  NOT_103(g8987,I14382);
  IV  NOT_104(g11546,g11519);
  IV  NOT_105(I10729,g5935);
  IV  NOT_106(g5253,g4346);
  IV  NOT_107(g7338,I11662);
  IV  NOT_108(I7509,g3566);
  IV  NOT_109(I9427,g4963);
  IV  NOT_110(g3800,g3292);
  IV  NOT_111(I15088,g9832);
  IV  NOT_112(g2907,I6074);
  IV  NOT_113(g7791,I12538);
  IV  NOT_114(I11143,g6446);
  IV  NOT_115(g6854,I10920);
  IV  NOT_116(g11088,I16871);
  IV  NOT_117(g7309,I11575);
  IV  NOT_118(g8299,I13255);
  IV  NOT_119(I9046,g4736);
  IV  NOT_120(g6941,g6503);
  IV  NOT_121(g2435,g201);
  IV  NOT_122(I14439,g8969);
  IV  NOT_123(g4010,g3144);
  IV  NOT_124(g2082,g1371);
  IV  NOT_125(I6932,g2850);
  IV  NOT_126(I7662,g3336);
  IV  NOT_127(I9446,g5052);
  IV  NOT_128(g5519,g4811);
  IV  NOT_129(g5740,I9302);
  IV  NOT_130(I5289,g49);
  IV  NOT_131(I9514,g5094);
  IV  NOT_132(g7808,I12589);
  IV  NOT_133(g2482,I5565);
  IV  NOT_134(I5658,g560);
  IV  NOT_135(I15497,g10119);
  IV  NOT_136(I6624,g2629);
  IV  NOT_137(g8892,I14242);
  IV  NOT_138(I11169,g6481);
  IV  NOT_139(g3213,I6388);
  IV  NOT_140(I6068,g2227);
  IV  NOT_141(g11497,I17510);
  IV  NOT_142(I13791,g8518);
  IV  NOT_143(I16867,g10913);
  IV  NOT_144(I10349,g6215);
  IV  NOT_145(g10260,g10125);
  IV  NOT_146(g7759,I12442);
  IV  NOT_147(I8473,g4577);
  IV  NOT_148(I14349,g8958);
  IV  NOT_149(g6708,I10689);
  IV  NOT_150(g10668,g10563);
  IV  NOT_151(I5271,g70);
  IV  NOT_152(I9191,g5546);
  IV  NOT_153(I9391,g5013);
  IV  NOT_154(g6219,g5426);
  IV  NOT_155(I15250,g9980);
  IV  NOT_156(I17100,g11221);
  IV  NOT_157(I14906,g9508);
  IV  NOT_158(g9825,I14976);
  IV  NOT_159(g7201,I11427);
  IV  NOT_160(I14083,g8747);
  IV  NOT_161(g10195,I15559);
  IV  NOT_162(I8324,g4794);
  IV  NOT_163(g6031,I9642);
  IV  NOT_164(g2915,I6094);
  IV  NOT_165(I13666,g8292);
  IV  NOT_166(I9695,g5212);
  IV  NOT_167(I11363,g6595);
  IV  NOT_168(I11217,g6529);
  IV  NOT_169(g6431,g6145);
  IV  NOT_170(g6252,I10015);
  IV  NOT_171(g4172,I7333);
  IV  NOT_172(g6812,I10846);
  IV  NOT_173(g8991,I14394);
  IV  NOT_174(g4372,I7677);
  IV  NOT_175(g7049,I11228);
  IV  NOT_176(I6576,g2617);
  IV  NOT_177(g10525,g10499);
  IV  NOT_178(g10488,I16101);
  IV  NOT_179(I10566,g5904);
  IV  NOT_180(I13478,g8191);
  IV  NOT_181(g5586,I8996);
  IV  NOT_182(g8709,g8674);
  IV  NOT_183(g2214,g115);
  IV  NOT_184(I9536,g5008);
  IV  NOT_185(g6176,I9905);
  IV  NOT_186(g4618,g3829);
  IV  NOT_187(I15296,g9995);
  IV  NOT_188(g4143,I7291);
  IV  NOT_189(I7381,g4078);
  IV  NOT_190(I9159,g5033);
  IV  NOT_191(g11339,I17142);
  IV  NOT_192(g8140,I13017);
  IV  NOT_193(I16979,g11088);
  IV  NOT_194(I16496,g10707);
  IV  NOT_195(g8078,I12936);
  IV  NOT_196(I7847,g3435);
  IV  NOT_197(I9359,g5576);
  IV  NOT_198(g8340,I13400);
  IV  NOT_199(g2110,I5002);
  IV  NOT_200(I15338,g10013);
  IV  NOT_201(g6405,g6133);
  IV  NOT_202(g8478,I13678);
  IV  NOT_203(I16111,g10385);
  IV  NOT_204(g4282,g4013);
  IV  NOT_205(g11644,I17736);
  IV  NOT_206(g7604,I12162);
  IV  NOT_207(g9768,g9432);
  IV  NOT_208(g4566,g3753);
  IV  NOT_209(g7098,I11333);
  IV  NOT_210(g10893,I16641);
  IV  NOT_211(I4961,g254);
  IV  NOT_212(g4988,I8358);
  IV  NOT_213(g6286,I10117);
  IV  NOT_214(g8959,I14326);
  IV  NOT_215(I13580,g8338);
  IV  NOT_216(I9016,g4722);
  IV  NOT_217(I6398,g2335);
  IV  NOT_218(g8517,I13720);
  IV  NOT_219(g3348,g2733);
  IV  NOT_220(I15060,g9696);
  IV  NOT_221(I15968,g10408);
  IV  NOT_222(I5332,g756);
  IV  NOT_223(g8482,g8329);
  IV  NOT_224(g2002,g818);
  IV  NOT_225(I10138,g5677);
  IV  NOT_226(g11060,g10937);
  IV  NOT_227(I17407,g11417);
  IV  NOT_228(I12303,g7242);
  IV  NOT_229(g5645,I9096);
  IV  NOT_230(I15855,g10336);
  IV  NOT_231(g2824,I5932);
  IV  NOT_232(g11197,g11112);
  IV  NOT_233(g4555,I7964);
  IV  NOT_234(g5691,g5236);
  IV  NOT_235(I9642,g5229);
  IV  NOT_236(g7539,I11953);
  IV  NOT_237(g7896,I12678);
  IV  NOT_238(g8656,I13941);
  IV  NOT_239(g9887,I15068);
  IV  NOT_240(I8199,g4013);
  IV  NOT_241(g6974,g6365);
  IV  NOT_242(g6270,I10069);
  IV  NOT_243(I14415,g8940);
  IV  NOT_244(g3260,I6428);
  IV  NOT_245(g11411,I17274);
  IV  NOT_246(I10852,g6751);
  IV  NOT_247(g10042,I15253);
  IV  NOT_248(g10255,g10139);
  IV  NOT_249(g6073,I9712);
  IV  NOT_250(g10189,I15545);
  IV  NOT_251(I4903,g259);
  IV  NOT_252(g2877,I6025);
  IV  NOT_253(I11531,g7126);
  IV  NOT_254(g10679,g10584);
  IV  NOT_255(g6796,g6252);
  IV  NOT_256(I8900,g4560);
  IV  NOT_257(I16735,g10855);
  IV  NOT_258(g1968,g369);
  IV  NOT_259(g5879,I9498);
  IV  NOT_260(I10963,g6793);
  IV  NOT_261(g10270,g10156);
  IV  NOT_262(g3463,g3256);
  IV  NOT_263(g7268,I11505);
  IV  NOT_264(g7362,I11734);
  IV  NOT_265(I11740,g7030);
  IV  NOT_266(g10188,I15542);
  IV  NOT_267(I12174,g6939);
  IV  NOT_268(I12796,g7543);
  IV  NOT_269(g5659,I9138);
  IV  NOT_270(g7419,g7206);
  IV  NOT_271(I15503,g10044);
  IV  NOT_272(I17441,g11445);
  IV  NOT_273(g6980,I11127);
  IV  NOT_274(I17206,g11323);
  IV  NOT_275(g4113,I7255);
  IV  NOT_276(g6069,I9706);
  IV  NOT_277(g11503,I17528);
  IV  NOT_278(g7052,I11235);
  IV  NOT_279(g8110,g7996);
  IV  NOT_280(g2556,g186);
  IV  NOT_281(g4313,g3586);
  IV  NOT_282(I16196,g10496);
  IV  NOT_283(I7817,g3399);
  IV  NOT_284(g8310,I13314);
  IV  NOT_285(g10460,I15971);
  IV  NOT_286(g2222,g158);
  IV  NOT_287(I11953,g6907);
  IV  NOT_288(I13373,g8226);
  IV  NOT_289(I6818,g2758);
  IV  NOT_290(g4202,I7423);
  IV  NOT_291(I6867,g2949);
  IV  NOT_292(I9880,g5405);
  IV  NOT_293(g10093,I15326);
  IV  NOT_294(I10484,g6155);
  IV  NOT_295(g9845,g9679);
  IV  NOT_296(g3720,I6888);
  IV  NOT_297(g10267,g10130);
  IV  NOT_298(g10294,I15704);
  IV  NOT_299(I11800,g7246);
  IV  NOT_300(g4908,g4396);
  IV  NOT_301(g5111,I8499);
  IV  NOT_302(g11450,I17407);
  IV  NOT_303(I13800,g8500);
  IV  NOT_304(g5275,g4371);
  IV  NOT_305(I11417,g6638);
  IV  NOT_306(I17758,g11647);
  IV  NOT_307(g3318,g2245);
  IV  NOT_308(g11315,I17108);
  IV  NOT_309(g4094,g2744);
  IV  NOT_310(I17435,g11454);
  IV  NOT_311(g10065,I15293);
  IV  NOT_312(I5092,g32);
  IV  NOT_313(g8002,I12832);
  IV  NOT_314(g5615,I9043);
  IV  NOT_315(g4567,g3374);
  IV  NOT_316(I8259,g4590);
  IV  NOT_317(g11202,g11112);
  IV  NOT_318(g7728,I12369);
  IV  NOT_319(g6287,I10120);
  IV  NOT_320(I14312,g8814);
  IV  NOT_321(I9612,g5149);
  IV  NOT_322(g10875,I16595);
  IV  NOT_323(I9243,g5245);
  IV  NOT_324(g11055,g10950);
  IV  NOT_325(g3393,g3144);
  IV  NOT_326(g9807,g9490);
  IV  NOT_327(g11111,g10974);
  IV  NOT_328(g4776,g3586);
  IV  NOT_329(I9935,g5477);
  IV  NOT_330(g4593,I8004);
  IV  NOT_331(I11964,g6910);
  IV  NOT_332(I7441,g3473);
  IV  NOT_333(I15986,g10417);
  IV  NOT_334(g3971,I7104);
  IV  NOT_335(g7070,I11289);
  IV  NOT_336(g2237,g713);
  IV  NOT_337(g6399,I10305);
  IV  NOT_338(g5284,g4376);
  IV  NOT_339(I11423,g6488);
  IV  NOT_340(g7470,g6927);
  IV  NOT_341(I15741,g10260);
  IV  NOT_342(g7897,g7712);
  IV  NOT_343(g7025,g6400);
  IV  NOT_344(I6370,g2356);
  IV  NOT_345(g7425,g7214);
  IV  NOT_346(I11587,g6828);
  IV  NOT_347(g2844,I5966);
  IV  NOT_348(I12553,g7676);
  IV  NOT_349(I12862,g7638);
  IV  NOT_350(I8215,g3981);
  IV  NOT_351(I10813,g6397);
  IV  NOT_352(g11384,I17209);
  IV  NOT_353(I14799,g9661);
  IV  NOT_354(I6821,g3015);
  IV  NOT_355(g2194,g47);
  IV  NOT_356(g10160,I15476);
  IV  NOT_357(g6797,I10801);
  IV  NOT_358(g11067,g10974);
  IV  NOT_359(g9342,I14531);
  IV  NOT_360(I12326,g7246);
  IV  NOT_361(g8928,I14257);
  IV  NOT_362(g3121,g2462);
  IV  NOT_363(I16280,g10537);
  IV  NOT_364(g4160,I7303);
  IV  NOT_365(g3321,I6484);
  IV  NOT_366(g2089,I4917);
  IV  NOT_367(g4933,I8298);
  IV  NOT_368(I14973,g9733);
  IV  NOT_369(g2731,I5789);
  IV  NOT_370(I16688,g10800);
  IV  NOT_371(I11543,g6881);
  IV  NOT_372(g5420,g4300);
  IV  NOT_373(I15801,g10282);
  IV  NOT_374(I12948,g8019);
  IV  NOT_375(g10455,I15956);
  IV  NOT_376(g8064,I12910);
  IV  NOT_377(g4521,g3586);
  IV  NOT_378(I14805,g9360);
  IV  NOT_379(g6291,I10132);
  IV  NOT_380(g2557,g1840);
  IV  NOT_381(g4050,I7163);
  IV  NOT_382(I13117,g7904);
  IV  NOT_383(I12904,g7985);
  IV  NOT_384(I4873,g105);
  IV  NOT_385(g8785,I14090);
  IV  NOT_386(g4450,g3914);
  IV  NOT_387(g5794,I9394);
  IV  NOT_388(g9097,g8892);
  IV  NOT_389(g2071,I4873);
  IV  NOT_390(g7678,I12307);
  IV  NOT_391(g6144,I9857);
  IV  NOT_392(I11569,g6821);
  IV  NOT_393(g3253,I6417);
  IV  NOT_394(I7743,g3762);
  IV  NOT_395(g6344,I10251);
  IV  NOT_396(g3938,g2991);
  IV  NOT_397(g7331,I11641);
  IV  NOT_398(I15196,g9974);
  IV  NOT_399(g9354,I14567);
  IV  NOT_400(g10201,g10175);
  IV  NOT_401(g7406,I11786);
  IV  NOT_402(g10277,I15675);
  IV  NOT_403(g2242,I5245);
  IV  NOT_404(I9213,g4944);
  IV  NOT_405(g3909,g2920);
  IV  NOT_406(I6106,g2116);
  IV  NOT_407(g7635,I12245);
  IV  NOT_408(I4869,g253);
  IV  NOT_409(I13568,g8343);
  IV  NOT_410(I13747,g8299);
  IV  NOT_411(I15526,g10051);
  IV  NOT_412(g8563,I13782);
  IV  NOT_413(g10075,I15302);
  IV  NOT_414(g4724,g3586);
  IV  NOT_415(g6259,I10036);
  IV  NOT_416(g4179,I7354);
  IV  NOT_417(g7766,I12463);
  IV  NOT_418(I5722,g2075);
  IV  NOT_419(g7682,g7148);
  IV  NOT_420(I13242,g8267);
  IV  NOT_421(I17500,g11478);
  IV  NOT_422(g6694,I10663);
  IV  NOT_423(g4379,g3698);
  IV  NOT_424(g3519,g3164);
  IV  NOT_425(g7801,I12568);
  IV  NOT_426(g7305,I11563);
  IV  NOT_427(I7411,g4140);
  IV  NOT_428(g8295,I13239);
  IV  NOT_429(g2955,I6156);
  IV  NOT_430(I8136,g4144);
  IV  NOT_431(g5628,I9062);
  IV  NOT_432(I6061,g2246);
  IV  NOT_433(I12183,g7007);
  IV  NOT_434(g6852,I10914);
  IV  NOT_435(I11814,g7196);
  IV  NOT_436(g5515,g4429);
  IV  NOT_437(I6461,g2261);
  IV  NOT_438(g5630,I9068);
  IV  NOT_439(I12397,g7284);
  IV  NOT_440(I4917,g584);
  IV  NOT_441(g2254,g131);
  IV  NOT_442(g2814,I5916);
  IV  NOT_443(g11402,I17249);
  IV  NOT_444(g4289,g4013);
  IV  NOT_445(g7748,I12409);
  IV  NOT_446(g4777,g3992);
  IV  NOT_447(I11807,g6854);
  IV  NOT_448(g11457,I17424);
  IV  NOT_449(I9090,g5567);
  IV  NOT_450(g4835,I8192);
  IV  NOT_451(I14400,g8891);
  IV  NOT_452(g2350,I5424);
  IV  NOT_453(g7755,I12430);
  IV  NOT_454(g9267,g8892);
  IV  NOT_455(g9312,I14509);
  IV  NOT_456(I13639,g8321);
  IV  NOT_457(g2038,g1776);
  IV  NOT_458(I8943,g4585);
  IV  NOT_459(I16763,g10890);
  IV  NOT_460(I12933,g7899);
  IV  NOT_461(g7226,I11464);
  IV  NOT_462(g8089,g7934);
  IV  NOT_463(g10352,I15820);
  IV  NOT_464(g2438,g243);
  IV  NOT_465(I11293,g6516);
  IV  NOT_466(I13230,g8244);
  IV  NOT_467(g2773,I5858);
  IV  NOT_468(g4271,g3971);
  IV  NOT_469(I6904,g2820);
  IV  NOT_470(I12508,g7731);
  IV  NOT_471(I11638,g6948);
  IV  NOT_472(I12634,g7727);
  IV  NOT_473(g10155,I15461);
  IV  NOT_474(I17613,g11550);
  IV  NOT_475(g10822,I16534);
  IV  NOT_476(I4786,g109);
  IV  NOT_477(I6046,g2218);
  IV  NOT_478(I9056,g4753);
  IV  NOT_479(g6951,I11097);
  IV  NOT_480(g10266,g10129);
  IV  NOT_481(I8228,g4468);
  IV  NOT_482(I14005,g8631);
  IV  NOT_483(g10170,g10118);
  IV  NOT_484(I8465,g4807);
  IV  NOT_485(I16660,g10793);
  IV  NOT_486(g7045,g6435);
  IV  NOT_487(I10538,g5910);
  IV  NOT_488(I8934,g4271);
  IV  NOT_489(I5424,g910);
  IV  NOT_490(I5795,g2462);
  IV  NOT_491(g7445,I11845);
  IV  NOT_492(g6114,I9795);
  IV  NOT_493(I5737,g2100);
  IV  NOT_494(I6403,g2337);
  IV  NOT_495(I5809,g2356);
  IV  NOT_496(g6314,I10201);
  IV  NOT_497(I7713,g3750);
  IV  NOT_498(g9761,g9454);
  IV  NOT_499(I11841,g7226);
  IV  NOT_500(I11992,g7058);
  IV  NOT_501(I11391,g6387);
  IV  NOT_502(I9851,g5405);
  IV  NOT_503(g2212,g686);
  IV  NOT_504(I13391,g8178);
  IV  NOT_505(g6870,I10952);
  IV  NOT_506(g4674,I8050);
  IV  NOT_507(g8948,I14299);
  IV  NOT_508(g3141,g2563);
  IV  NOT_509(I6391,g2478);
  IV  NOT_510(I5672,g569);
  IV  NOT_511(I15688,g10207);
  IV  NOT_512(g5040,I8421);
  IV  NOT_513(I5077,g35);
  IV  NOT_514(g1983,g750);
  IV  NOT_515(g6825,I10873);
  IV  NOT_516(g3710,g3215);
  IV  NOT_517(g7369,g7273);
  IV  NOT_518(g7602,I12156);
  IV  NOT_519(g10167,I15497);
  IV  NOT_520(g10194,g10062);
  IV  NOT_521(g10589,I16252);
  IV  NOT_522(I16550,g10726);
  IV  NOT_523(g4541,I7946);
  IV  NOT_524(g7007,I11146);
  IV  NOT_525(I17371,g11410);
  IV  NOT_526(I17234,g11353);
  IV  NOT_527(g7920,g7516);
  IV  NOT_528(I11578,g6824);
  IV  NOT_529(I12574,g7522);
  IV  NOT_530(g10524,g10458);
  IV  NOT_531(g2229,g162);
  IV  NOT_532(I15157,g9931);
  IV  NOT_533(I16307,g10589);
  IV  NOT_534(g4332,g4130);
  IV  NOT_535(I12205,g6993);
  IV  NOT_536(g7767,I12466);
  IV  NOT_537(I6159,g2123);
  IV  NOT_538(g11157,g10950);
  IV  NOT_539(g4680,g3829);
  IV  NOT_540(g6136,I9845);
  IV  NOT_541(g8150,I13039);
  IV  NOT_542(g4209,I7444);
  IV  NOT_543(g4353,I7636);
  IV  NOT_544(g5666,I9159);
  IV  NOT_545(g6336,I10231);
  IV  NOT_546(g8350,I13430);
  IV  NOT_547(I13586,g8356);
  IV  NOT_548(g10119,I15365);
  IV  NOT_549(I8337,g4352);
  IV  NOT_550(g8438,I13612);
  IV  NOT_551(g6594,I10560);
  IV  NOT_552(g11066,g10974);
  IV  NOT_553(g4802,g3337);
  IV  NOT_554(I13442,g8182);
  IV  NOT_555(g8009,I12849);
  IV  NOT_556(I5304,g79);
  IV  NOT_557(g10118,I15362);
  IV  NOT_558(I6016,g2201);
  IV  NOT_559(I6757,g2732);
  IV  NOT_560(g7793,I12544);
  IV  NOT_561(I9279,g5314);
  IV  NOT_562(g5648,I9105);
  IV  NOT_563(g6806,I10828);
  IV  NOT_564(g5875,g5361);
  IV  NOT_565(g6943,I11079);
  IV  NOT_566(I16269,g10558);
  IV  NOT_567(I9720,g5248);
  IV  NOT_568(I12592,g7445);
  IV  NOT_569(g10616,I16289);
  IV  NOT_570(g4558,g3880);
  IV  NOT_571(g5655,I9126);
  IV  NOT_572(I13615,g8333);
  IV  NOT_573(g7415,I11797);
  IV  NOT_574(g7227,I11467);
  IV  NOT_575(I9872,g5557);
  IV  NOT_576(g10313,I15741);
  IV  NOT_577(I5926,g2172);
  IV  NOT_578(I13720,g8358);
  IV  NOT_579(I9652,g5426);
  IV  NOT_580(I5754,g2304);
  IV  NOT_581(I10991,g6759);
  IV  NOT_582(I15763,g10244);
  IV  NOT_583(I11275,g6502);
  IV  NOT_584(g10276,I15672);
  IV  NOT_585(g11511,I17552);
  IV  NOT_586(g4901,I8268);
  IV  NOT_587(I7760,g3768);
  IV  NOT_588(I16670,g10797);
  IV  NOT_589(I11746,g6857);
  IV  NOT_590(I13430,g8241);
  IV  NOT_591(g10305,I15725);
  IV  NOT_592(g10254,g10196);
  IV  NOT_593(g4511,g3586);
  IV  NOT_594(g10900,I16656);
  IV  NOT_595(g9576,I14713);
  IV  NOT_596(g2837,g2130);
  IV  NOT_597(g10466,I15989);
  IV  NOT_598(g5884,I9505);
  IV  NOT_599(I5044,g1182);
  IV  NOT_600(g6433,I10349);
  IV  NOT_601(g5839,I9452);
  IV  NOT_602(g8229,g7826);
  IV  NOT_603(I6654,g2952);
  IV  NOT_604(g8993,I14400);
  IV  NOT_605(g2620,g1998);
  IV  NOT_606(I12846,g7685);
  IV  NOT_607(g2462,I5555);
  IV  NOT_608(g9349,I14552);
  IV  NOT_609(I8815,g4471);
  IV  NOT_610(g10101,I15335);
  IV  NOT_611(g10177,I15523);
  IV  NOT_612(I16667,g10780);
  IV  NOT_613(I13806,g8478);
  IV  NOT_614(I7220,g3213);
  IV  NOT_615(I5862,g2537);
  IV  NOT_616(I9598,g5120);
  IV  NOT_617(I7779,g3774);
  IV  NOT_618(I17724,g11625);
  IV  NOT_619(g6845,I10907);
  IV  NOT_620(g7502,I11882);
  IV  NOT_621(I8154,g3636);
  IV  NOT_622(I10584,g5864);
  IV  NOT_623(I17359,g11372);
  IV  NOT_624(g3545,I6733);
  IV  NOT_625(I15314,g10007);
  IV  NOT_626(g11550,I17591);
  IV  NOT_627(I15287,g9980);
  IV  NOT_628(g6195,g5426);
  IV  NOT_629(I7423,g3331);
  IV  NOT_630(g6137,I9848);
  IV  NOT_631(g5667,I9162);
  IV  NOT_632(g6395,I10293);
  IV  NOT_633(g3380,I6576);
  IV  NOT_634(g5143,g4682);
  IV  NOT_635(g6337,I10234);
  IV  NOT_636(I16487,g10771);
  IV  NOT_637(g6913,I11021);
  IV  NOT_638(g10064,I15290);
  IV  NOT_639(g11287,g11207);
  IV  NOT_640(I15085,g9720);
  IV  NOT_641(g2249,g127);
  IV  NOT_642(I9625,g5405);
  IV  NOT_643(g4580,g3880);
  IV  NOT_644(I10759,g5803);
  IV  NOT_645(g11307,I17092);
  IV  NOT_646(g11076,I16843);
  IV  NOT_647(I9232,g4944);
  IV  NOT_648(g7188,I11408);
  IV  NOT_649(g7689,I12322);
  IV  NOT_650(I17121,g11231);
  IV  NOT_651(g11596,g11580);
  IV  NOT_652(g7388,I11773);
  IV  NOT_653(I10114,g5768);
  IV  NOT_654(I9253,g5052);
  IV  NOT_655(I9938,g5478);
  IV  NOT_656(g10874,I16592);
  IV  NOT_657(g11054,g10950);
  IV  NOT_658(g6807,I10831);
  IV  NOT_659(I9813,g5241);
  IV  NOT_660(I6417,g2344);
  IV  NOT_661(g5693,I9224);
  IV  NOT_662(g11243,g11112);
  IV  NOT_663(I17344,g11369);
  IV  NOT_664(g3507,g3307);
  IV  NOT_665(g4262,g4013);
  IV  NOT_666(g2298,I5336);
  IV  NOT_667(g2085,I4903);
  IV  NOT_668(I7665,g3732);
  IV  NOT_669(g10630,I16311);
  IV  NOT_670(g11431,I17344);
  IV  NOT_671(g6859,I10937);
  IV  NOT_672(g7028,g6407);
  IV  NOT_673(I6982,g2889);
  IV  NOT_674(g6266,I10057);
  IV  NOT_675(I15269,g9993);
  IV  NOT_676(g10166,I15494);
  IV  NOT_677(g7030,I11183);
  IV  NOT_678(I12583,g7546);
  IV  NOT_679(I9519,g4998);
  IV  NOT_680(g8062,I12904);
  IV  NOT_681(g7430,g7221);
  IV  NOT_682(I15341,g10019);
  IV  NOT_683(I5414,g904);
  IV  NOT_684(I16286,g10540);
  IV  NOT_685(I7999,g4114);
  IV  NOT_686(g2854,I5986);
  IV  NOT_687(I17173,g11293);
  IV  NOT_688(I5946,g2176);
  IV  NOT_689(I10849,g6734);
  IV  NOT_690(g11341,I17146);
  IV  NOT_691(I7633,g3474);
  IV  NOT_692(g4889,I8240);
  IV  NOT_693(g2941,I6118);
  IV  NOT_694(g6248,I10003);
  IV  NOT_695(g11655,I17767);
  IV  NOT_696(g9258,g8892);
  IV  NOT_697(g3905,g2920);
  IV  NOT_698(g10892,I16638);
  IV  NOT_699(g9818,I14955);
  IV  NOT_700(g9352,I14561);
  IV  NOT_701(I7303,g3262);
  IV  NOT_702(I8293,g4779);
  IV  NOT_703(I10398,g5820);
  IV  NOT_704(I13475,g8173);
  IV  NOT_705(g11180,I16941);
  IV  NOT_706(g7826,I12627);
  IV  NOT_707(g3628,g3111);
  IV  NOT_708(g6255,I10024);
  IV  NOT_709(g4175,I7342);
  IV  NOT_710(g6081,g4977);
  IV  NOT_711(g6815,I10855);
  IV  NOT_712(I10141,g5683);
  IV  NOT_713(g4375,g3638);
  IV  NOT_714(I10804,g6388);
  IV  NOT_715(I5513,g255);
  IV  NOT_716(g3630,I6789);
  IV  NOT_717(g8788,I14097);
  IV  NOT_718(I11222,g6533);
  IV  NOT_719(I12282,g7113);
  IV  NOT_720(I15335,g10007);
  IV  NOT_721(I16601,g10806);
  IV  NOT_722(g5113,I8503);
  IV  NOT_723(g6692,I10659);
  IV  NOT_724(I16187,g10492);
  IV  NOT_725(g6097,I9754);
  IV  NOT_726(I7732,g3758);
  IV  NOT_727(g7910,g7460);
  IV  NOT_728(I12357,g7147);
  IV  NOT_729(g2219,g94);
  IV  NOT_730(g9893,I15082);
  IV  NOT_731(g2640,g1984);
  IV  NOT_732(g6154,I9875);
  IV  NOT_733(g4285,g3688);
  IV  NOT_734(g6354,g5867);
  IV  NOT_735(g2031,g1690);
  IV  NOT_736(g10907,I16673);
  IV  NOT_737(g5202,g4640);
  IV  NOT_738(g6960,I11112);
  IV  NOT_739(I15694,g10234);
  IV  NOT_740(I5378,g1857);
  IV  NOT_741(g2431,I5510);
  IV  NOT_742(I15965,g10405);
  IV  NOT_743(g2252,I5271);
  IV  NOT_744(g2812,g2158);
  IV  NOT_745(I7240,g2824);
  IV  NOT_746(g7609,I12177);
  IV  NOT_747(I10135,g6249);
  IV  NOT_748(g7308,I11572);
  IV  NOT_749(g8192,I13117);
  IV  NOT_750(g2958,I6163);
  IV  NOT_751(g8085,g7932);
  IV  NOT_752(g10074,I15299);
  IV  NOT_753(g5094,I8462);
  IV  NOT_754(I13347,g8122);
  IV  NOT_755(g2176,g82);
  IV  NOT_756(g9026,I14415);
  IV  NOT_757(g8485,g8341);
  IV  NOT_758(g4184,I7369);
  IV  NOT_759(g5494,g4412);
  IV  NOT_760(g3750,I6941);
  IV  NOT_761(g2005,g928);
  IV  NOT_762(g7883,g7689);
  IV  NOT_763(I7043,g2908);
  IV  NOT_764(g4384,I7707);
  IV  NOT_765(I9141,g5402);
  IV  NOT_766(I9860,g5405);
  IV  NOT_767(g5567,I8982);
  IV  NOT_768(g4339,g4144);
  IV  NOT_769(I9341,g5013);
  IV  NOT_770(g10238,g10191);
  IV  NOT_771(I16169,g10448);
  IV  NOT_772(I9525,g5001);
  IV  NOT_773(I14361,g8951);
  IV  NOT_774(g2829,I5943);
  IV  NOT_775(g11619,I17675);
  IV  NOT_776(g2765,g2184);
  IV  NOT_777(g9821,I14964);
  IV  NOT_778(g11502,I17525);
  IV  NOT_779(g7758,I12439);
  IV  NOT_780(I5916,g2217);
  IV  NOT_781(I13236,g8245);
  IV  NOT_782(g7066,I11275);
  IV  NOT_783(g7589,I12099);
  IV  NOT_784(g4424,g3688);
  IV  NOT_785(g3040,g2135);
  IV  NOT_786(g4737,g3440);
  IV  NOT_787(I11351,g6698);
  IV  NOT_788(I13952,g8451);
  IV  NOT_789(g5593,I9013);
  IV  NOT_790(g6112,I9789);
  IV  NOT_791(I13351,g8214);
  IV  NOT_792(g6218,I9965);
  IV  NOT_793(g6267,I10060);
  IV  NOT_794(g3440,g3041);
  IV  NOT_795(g6312,I10195);
  IV  NOT_796(g11618,I17672);
  IV  NOT_797(g9984,I15184);
  IV  NOT_798(I11821,g7205);
  IV  NOT_799(g10176,I15520);
  IV  NOT_800(g10185,g10040);
  IV  NOT_801(g10675,g10574);
  IV  NOT_802(I16479,g10767);
  IV  NOT_803(g10092,I15323);
  IV  NOT_804(I10048,g5734);
  IV  NOT_805(I16363,g10599);
  IV  NOT_806(I16217,g10501);
  IV  NOT_807(g3323,g2157);
  IV  NOT_808(I15278,g10033);
  IV  NOT_809(g7571,I12035);
  IV  NOT_810(g7365,I11743);
  IV  NOT_811(g2733,I5795);
  IV  NOT_812(g4077,I7202);
  IV  NOT_813(g6001,I9625);
  IV  NOT_814(g7048,I11225);
  IV  NOT_815(g10154,I15458);
  IV  NOT_816(g2270,I5311);
  IV  NOT_817(I5798,g2085);
  IV  NOT_818(I17240,g11395);
  IV  NOT_819(g7711,I12344);
  IV  NOT_820(g4523,g3546);
  IV  NOT_821(I10221,g6117);
  IV  NOT_822(I11790,g7246);
  IV  NOT_823(g8520,I13729);
  IV  NOT_824(g6293,I10138);
  IV  NOT_825(g11469,I17444);
  IV  NOT_826(g8219,g7826);
  IV  NOT_827(g2225,I5210);
  IV  NOT_828(g8640,g8512);
  IV  NOT_829(g10935,g10827);
  IV  NOT_830(g2610,I5731);
  IV  NOT_831(g2073,I4879);
  IV  NOT_832(g2796,g2276);
  IV  NOT_833(g11468,I17441);
  IV  NOT_834(g11039,I16778);
  IV  NOT_835(I6851,g2937);
  IV  NOT_836(g4205,I7432);
  IV  NOT_837(I7697,g3743);
  IV  NOT_838(I10613,g6000);
  IV  NOT_839(I11873,g6863);
  IV  NOT_840(g10883,g10809);
  IV  NOT_841(I17755,g11646);
  IV  NOT_842(g7333,I11647);
  IV  NOT_843(g9106,I14439);
  IV  NOT_844(I7210,g2798);
  IV  NOT_845(g7774,I12487);
  IV  NOT_846(g5521,g4530);
  IV  NOT_847(g3528,g3164);
  IV  NOT_848(g8958,I14323);
  IV  NOT_849(I16580,g10826);
  IV  NOT_850(I17770,g11649);
  IV  NOT_851(g11038,I16775);
  IV  NOT_852(g5050,I8429);
  IV  NOT_853(g2124,I5050);
  IV  NOT_854(g3351,I6535);
  IV  NOT_855(g5641,I9084);
  IV  NOT_856(I17563,g11492);
  IV  NOT_857(g2980,g1983);
  IV  NOT_858(g6727,g5997);
  IV  NOT_859(g8376,I13478);
  IV  NOT_860(I5632,g932);
  IV  NOT_861(I5095,g37);
  IV  NOT_862(I6260,g2025);
  IV  NOT_863(g2069,I4869);
  IV  NOT_864(I9111,g5596);
  IV  NOT_865(g7196,I11420);
  IV  NOT_866(g4551,g3946);
  IV  NOT_867(I15601,g10173);
  IV  NOT_868(I9311,g4915);
  IV  NOT_869(I15187,g9968);
  IV  NOT_870(g7803,I12574);
  IV  NOT_871(I12248,g7098);
  IV  NOT_872(I13209,g8198);
  IV  NOT_873(g4499,g3546);
  IV  NOT_874(I8848,g4490);
  IV  NOT_875(g2540,I5655);
  IV  NOT_876(g7538,I11950);
  IV  NOT_877(I13834,g8488);
  IV  NOT_878(I5579,g1197);
  IV  NOT_879(g7780,I12505);
  IV  NOT_880(g5724,I9268);
  IV  NOT_881(g9027,I14418);
  IV  NOT_882(g2206,I5171);
  IV  NOT_883(I12779,g7608);
  IV  NOT_884(g10729,g10630);
  IV  NOT_885(g6703,I10678);
  IV  NOT_886(I9174,g4903);
  IV  NOT_887(I5719,g2072);
  IV  NOT_888(g10577,g10526);
  IV  NOT_889(I17767,g11648);
  IV  NOT_890(g7509,I11889);
  IV  NOT_891(g9427,g9079);
  IV  NOT_892(I10033,g5693);
  IV  NOT_893(I7820,g3811);
  IV  NOT_894(I10234,g6114);
  IV  NOT_895(g4754,g3440);
  IV  NOT_896(I16531,g10720);
  IV  NOT_897(g10439,g10334);
  IV  NOT_898(I11021,g6398);
  IV  NOT_899(I12081,g6934);
  IV  NOT_900(g5878,g5309);
  IV  NOT_901(g6932,I11058);
  IV  NOT_902(g7662,I12279);
  IV  NOT_903(g4273,g4013);
  IV  NOT_904(I16178,g10490);
  IV  NOT_905(I12786,g7622);
  IV  NOT_906(I17633,g11578);
  IV  NOT_907(g5658,I9135);
  IV  NOT_908(g5777,I9365);
  IV  NOT_909(I10795,g6123);
  IV  NOT_910(I13726,g8375);
  IV  NOT_911(g7467,g7148);
  IV  NOT_912(g1990,g774);
  IV  NOT_913(I6118,g2248);
  IV  NOT_914(g8225,g7826);
  IV  NOT_915(I17191,g11315);
  IV  NOT_916(I17719,g11623);
  IV  NOT_917(I11614,g6838);
  IV  NOT_918(g8610,g8483);
  IV  NOT_919(I6367,g2045);
  IV  NOT_920(I9180,g4905);
  IV  NOT_921(I12647,g7711);
  IV  NOT_922(I16676,g10798);
  IV  NOT_923(I16685,g10785);
  IV  NOT_924(I11436,g6488);
  IV  NOT_925(I9380,g5013);
  IV  NOT_926(g10349,I15811);
  IV  NOT_927(g9345,I14540);
  IV  NOT_928(I16953,g11082);
  IV  NOT_929(I13436,g8187);
  IV  NOT_930(I9591,g5095);
  IV  NOT_931(I16373,g10593);
  IV  NOT_932(g4444,I7800);
  IV  NOT_933(g8473,I13669);
  IV  NOT_934(g2199,g48);
  IV  NOT_935(g11410,I17271);
  IV  NOT_936(g2399,g605);
  IV  NOT_937(g9763,I14906);
  IV  NOT_938(g7093,I11326);
  IV  NOT_939(I12999,g7844);
  IV  NOT_940(g3372,g3121);
  IV  NOT_941(I10514,g6154);
  IV  NOT_942(I12380,g7204);
  IV  NOT_943(g10906,I16670);
  IV  NOT_944(I15479,g10091);
  IV  NOT_945(I13320,g8096);
  IV  NOT_946(g10083,I15311);
  IV  NOT_947(I9020,g4773);
  IV  NOT_948(g8124,g8011);
  IV  NOT_949(g10284,g10167);
  IV  NOT_950(g7256,I11489);
  IV  NOT_951(g8980,I14361);
  IV  NOT_952(g7816,I12613);
  IV  NOT_953(g8324,I13354);
  IV  NOT_954(g11479,I17470);
  IV  NOT_955(I6193,g2155);
  IV  NOT_956(I11593,g6830);
  IV  NOT_957(g3143,I6363);
  IV  NOT_958(g11363,I17188);
  IV  NOT_959(g3343,g2779);
  IV  NOT_960(I11122,g6450);
  IV  NOT_961(g2797,g2524);
  IV  NOT_962(I13122,g7966);
  IV  NOT_963(I6549,g2838);
  IV  NOT_964(g4543,g3946);
  IV  NOT_965(I10421,g5826);
  IV  NOT_966(I11464,g6443);
  IV  NOT_967(g3566,I6738);
  IV  NOT_968(I6971,g2882);
  IV  NOT_969(g6716,g5949);
  IV  NOT_970(I14421,g8944);
  IV  NOT_971(g2245,I5254);
  IV  NOT_972(g6149,I9866);
  IV  NOT_973(g3988,g3121);
  IV  NOT_974(I6686,g3015);
  IV  NOT_975(g6349,I10258);
  IV  NOT_976(g7847,I12638);
  IV  NOT_977(g3693,g2920);
  IV  NOT_978(I11034,g6629);
  IV  NOT_979(I10012,g5543);
  IV  NOT_980(g3334,I6517);
  IV  NOT_981(I5725,g2079);
  IV  NOT_982(g7685,g7148);
  IV  NOT_983(g7197,I11423);
  IV  NOT_984(I11641,g6960);
  IV  NOT_985(I11797,g6852);
  IV  NOT_986(g5997,I9617);
  IV  NOT_987(I15580,g10155);
  IV  NOT_988(I13797,g8473);
  IV  NOT_989(I6598,g2623);
  IV  NOT_990(g7021,I11162);
  IV  NOT_991(g4729,g3586);
  IV  NOT_992(g4961,I8333);
  IV  NOT_993(g7421,I11807);
  IV  NOT_994(g10139,I15415);
  IV  NOT_995(g2344,I5410);
  IV  NOT_996(I8211,g3566);
  IV  NOT_997(I9905,g5300);
  IV  NOT_998(g6398,I10302);
  IV  NOT_999(I10541,g6176);
  IV  NOT_1000(I6121,g2121);
  IV  NOT_1001(g1963,g110);
  IV  NOT_1002(I17324,g11347);
  IV  NOT_1003(g7263,I11498);
  IV  NOT_1004(I14473,g8921);
  IV  NOT_1005(g2207,I5174);
  IV  NOT_1006(g10138,I15412);
  IV  NOT_1007(I17701,g11617);
  IV  NOT_1008(I10789,g5867);
  IV  NOT_1009(I12448,g7530);
  IV  NOT_1010(I13409,g8141);
  IV  NOT_1011(I17534,g11495);
  IV  NOT_1012(g3792,I7017);
  IV  NOT_1013(g5353,I8820);
  IV  NOT_1014(g8849,g8745);
  IV  NOT_1015(g2259,I5292);
  IV  NOT_1016(g6241,I9992);
  IV  NOT_1017(g2819,g2159);
  IV  NOT_1018(I11408,g6405);
  IV  NOT_1019(I12505,g7728);
  IV  NOT_1020(I11635,g6947);
  IV  NOT_1021(I10724,g6096);
  IV  NOT_1022(g11084,I16863);
  IV  NOT_1023(g4885,I8228);
  IV  NOT_1024(g4414,I7752);
  IV  NOT_1025(I10325,g6003);
  IV  NOT_1026(g11110,g10974);
  IV  NOT_1027(g3621,I6754);
  IV  NOT_1028(I6938,g2854);
  IV  NOT_1029(I7668,g3733);
  IV  NOT_1030(g2852,I5982);
  IV  NOT_1031(I7840,g3431);
  IV  NOT_1032(I16543,g10747);
  IV  NOT_1033(g10852,g10740);
  IV  NOT_1034(g8781,I14080);
  IV  NOT_1035(I8614,g4414);
  IV  NOT_1036(I10920,g6733);
  IV  NOT_1037(I10535,g5867);
  IV  NOT_1038(I12026,g7119);
  IV  NOT_1039(I10434,g5843);
  IV  NOT_1040(g11179,I16938);
  IV  NOT_1041(g2701,g2040);
  IV  NOT_1042(g3113,I6343);
  IV  NOT_1043(g7562,g6984);
  IV  NOT_1044(I14358,g8950);
  IV  NOT_1045(I7390,g4087);
  IV  NOT_1046(I10828,g6708);
  IV  NOT_1047(I10946,g6548);
  IV  NOT_1048(g8797,I14116);
  IV  NOT_1049(g6644,I10601);
  IV  NOT_1050(g4513,g3546);
  IV  NOT_1051(g7631,I12235);
  IV  NOT_1052(I5171,g1419);
  IV  NOT_1053(g7723,I12354);
  IV  NOT_1054(g6119,I9810);
  IV  NOT_1055(I9973,g5502);
  IV  NOT_1056(g7817,I12616);
  IV  NOT_1057(g5901,g5361);
  IV  NOT_1058(I4920,g260);
  IV  NOT_1059(g8291,I13227);
  IV  NOT_1060(g11373,I17198);
  IV  NOT_1061(g3094,I6302);
  IV  NOT_1062(g6258,I10033);
  IV  NOT_1063(g4178,I7351);
  IV  NOT_1064(g4436,g3638);
  IV  NOT_1065(g6818,I10864);
  IV  NOT_1066(g4679,g4013);
  IV  NOT_1067(g11654,I17764);
  IV  NOT_1068(g4378,I7697);
  IV  NOT_1069(g7605,I12165);
  IV  NOT_1070(g5511,I8934);
  IV  NOT_1071(I11575,g6823);
  IV  NOT_1072(g3518,g3164);
  IV  NOT_1073(I10682,g6051);
  IV  NOT_1074(g10576,g10524);
  IV  NOT_1075(I9040,g4794);
  IV  NOT_1076(g8144,I13027);
  IV  NOT_1077(g8344,I13412);
  IV  NOT_1078(g6717,I10706);
  IV  NOT_1079(I9440,g5078);
  IV  NOT_1080(g11417,I17302);
  IV  NOT_1081(I13711,g8342);
  IV  NOT_1082(I16814,g10910);
  IV  NOT_1083(I12433,g7657);
  IV  NOT_1084(g4335,I7612);
  IV  NOT_1085(I9123,g4890);
  IV  NOT_1086(I11109,g6464);
  IV  NOT_1087(g7751,I12418);
  IV  NOT_1088(g4182,I7363);
  IV  NOT_1089(I9323,g5620);
  IV  NOT_1090(I13109,g7981);
  IV  NOT_1091(g4288,g4130);
  IV  NOT_1092(I11537,g7144);
  IV  NOT_1093(g4382,g3638);
  IV  NOT_1094(I16772,g10887);
  IV  NOT_1095(g3776,g2579);
  IV  NOT_1096(g6893,I10991);
  IV  NOT_1097(g5574,g4300);
  IV  NOT_1098(g5864,I9483);
  IV  NOT_1099(g10200,g10169);
  IV  NOT_1100(g8694,I13975);
  IV  NOT_1101(g2825,I5935);
  IV  NOT_1102(g2650,g2006);
  IV  NOT_1103(g10608,I16283);
  IV  NOT_1104(g10115,I15353);
  IV  NOT_1105(g6386,I10282);
  IV  NOT_1106(g7585,I12081);
  IV  NOT_1107(I17447,g11457);
  IV  NOT_1108(I5684,g572);
  IV  NOT_1109(I8061,g3381);
  IV  NOT_1110(g4805,g3337);
  IV  NOT_1111(I7163,g2643);
  IV  NOT_1112(I5963,g2179);
  IV  NOT_1113(I7810,g3799);
  IV  NOT_1114(g7041,g6427);
  IV  NOT_1115(I7363,g4005);
  IV  NOT_1116(I16638,g10863);
  IV  NOT_1117(g2008,g971);
  IV  NOT_1118(I13606,g8311);
  IV  NOT_1119(I12971,g8039);
  IV  NOT_1120(I11303,g6526);
  IV  NOT_1121(g6274,I10081);
  IV  NOT_1122(I7432,g3663);
  IV  NOT_1123(g6426,I10340);
  IV  NOT_1124(g11423,I17324);
  IV  NOT_1125(g2336,g1900);
  IV  NOT_1126(I16416,g10664);
  IV  NOT_1127(I12369,g7189);
  IV  NOT_1128(I9875,g5278);
  IV  NOT_1129(I7453,g3708);
  IV  NOT_1130(g6170,g5426);
  IV  NOT_1131(I14506,g8923);
  IV  NOT_1132(g7673,I12296);
  IV  NOT_1133(I9655,g5173);
  IV  NOT_1134(g6125,I9822);
  IV  NOT_1135(I5707,g2418);
  IV  NOT_1136(g8886,I14228);
  IV  NOT_1137(g3521,g3164);
  IV  NOT_1138(g8951,I14306);
  IV  NOT_1139(I16510,g10712);
  IV  NOT_1140(g5262,g4353);
  IV  NOT_1141(g3050,I6260);
  IV  NOT_1142(I11091,g6657);
  IV  NOT_1143(g10973,I16720);
  IV  NOT_1144(g5736,I9296);
  IV  NOT_1145(g6984,g6382);
  IV  NOT_1146(g6280,I10099);
  IV  NOT_1147(g6939,I11071);
  IV  NOT_1148(g7669,I12286);
  IV  NOT_1149(I17246,g11341);
  IV  NOT_1150(g11543,g11519);
  IV  NOT_1151(g3996,g3144);
  IV  NOT_1152(g10184,g10039);
  IV  NOT_1153(I12412,g7520);
  IV  NOT_1154(I8403,g4264);
  IV  NOT_1155(g10674,g10584);
  IV  NOT_1156(g8314,I13326);
  IV  NOT_1157(g5623,I9053);
  IV  NOT_1158(g7772,I12481);
  IV  NOT_1159(I7157,g3015);
  IV  NOT_1160(g7058,I11255);
  IV  NOT_1161(I12133,g6870);
  IV  NOT_1162(I5957,g2178);
  IV  NOT_1163(I7357,g4077);
  IV  NOT_1164(g2122,I5044);
  IV  NOT_1165(g2228,g28);
  IV  NOT_1166(g7531,I11929);
  IV  NOT_1167(g4095,I7233);
  IV  NOT_1168(g9554,I14697);
  IV  NOT_1169(g8870,I14182);
  IV  NOT_1170(g2322,I5378);
  IV  NOT_1171(I10927,g6755);
  IV  NOT_1172(g7458,g7123);
  IV  NOT_1173(g5889,I9514);
  IV  NOT_1174(I12229,g7070);
  IV  NOT_1175(I6962,g2791);
  IV  NOT_1176(g4495,I7886);
  IV  NOT_1177(I9839,g5226);
  IV  NOT_1178(g2230,g704);
  IV  NOT_1179(g4437,g3345);
  IV  NOT_1180(g4102,I7244);
  IV  NOT_1181(I17591,g11514);
  IV  NOT_1182(g4208,I7441);
  IV  NOT_1183(g7890,g7479);
  IV  NOT_1184(g8650,I13933);
  IV  NOT_1185(I13840,g8488);
  IV  NOT_1186(I16586,g10850);
  IV  NOT_1187(g3379,g3121);
  IV  NOT_1188(I15568,g10094);
  IV  NOT_1189(g10934,g10827);
  IV  NOT_1190(g6106,I9773);
  IV  NOT_1191(g5175,g4682);
  IV  NOT_1192(g6306,I10177);
  IV  NOT_1193(g7505,g7148);
  IV  NOT_1194(g3878,g2920);
  IV  NOT_1195(g11242,g11112);
  IV  NOT_1196(I5098,g38);
  IV  NOT_1197(g8008,I12846);
  IV  NOT_1198(I10240,g5937);
  IV  NOT_1199(g7011,g6503);
  IV  NOT_1200(g4719,g3586);
  IV  NOT_1201(g10692,I16363);
  IV  NOT_1202(g5651,I9114);
  IV  NOT_1203(I6587,g2620);
  IV  NOT_1204(I10648,g6030);
  IV  NOT_1205(I15814,g10202);
  IV  NOT_1206(g8336,I13388);
  IV  NOT_1207(I14903,g9507);
  IV  NOT_1208(I5833,g2103);
  IV  NOT_1209(g6387,g6121);
  IV  NOT_1210(g5285,g4355);
  IV  NOT_1211(g6461,I10391);
  IV  NOT_1212(I15807,g10284);
  IV  NOT_1213(I15974,g10411);
  IV  NOT_1214(I8858,g4506);
  IV  NOT_1215(g2550,g1834);
  IV  NOT_1216(g7074,I11299);
  IV  NOT_1217(I16720,g10854);
  IV  NOT_1218(g3271,I6443);
  IV  NOT_1219(g10400,g10348);
  IV  NOT_1220(g2845,g2168);
  IV  NOT_1221(I9282,g5633);
  IV  NOT_1222(I15639,g10179);
  IV  NOT_1223(I10563,g6043);
  IV  NOT_1224(I5584,g1200);
  IV  NOT_1225(g10214,I15586);
  IV  NOT_1226(g9490,g9324);
  IV  NOT_1227(g9823,I14970);
  IV  NOT_1228(g2195,g83);
  IV  NOT_1229(g4265,g3664);
  IV  NOT_1230(I15293,g10001);
  IV  NOT_1231(I9988,g5526);
  IV  NOT_1232(g6427,I10343);
  IV  NOT_1233(I12627,g7697);
  IV  NOT_1234(g2395,g231);
  IV  NOT_1235(g2891,I6055);
  IV  NOT_1236(g5184,g4682);
  IV  NOT_1237(g2337,I5395);
  IV  NOT_1238(I11483,g6567);
  IV  NOT_1239(g2913,I6088);
  IV  NOT_1240(g10329,I15775);
  IV  NOT_1241(g10207,g10186);
  IV  NOT_1242(g4442,g3638);
  IV  NOT_1243(I6985,g2890);
  IV  NOT_1244(g6904,I11008);
  IV  NOT_1245(g6200,I9935);
  IV  NOT_1246(g11638,I17724);
  IV  NOT_1247(g10539,I16184);
  IV  NOT_1248(g4786,I8154);
  IV  NOT_1249(g6046,I9669);
  IV  NOT_1250(g8065,I12913);
  IV  NOT_1251(g3799,I7022);
  IV  NOT_1252(I8315,g4788);
  IV  NOT_1253(I8811,g4465);
  IV  NOT_1254(g6446,I10370);
  IV  NOT_1255(g8122,I12981);
  IV  NOT_1256(g3981,I7118);
  IV  NOT_1257(g8465,g8289);
  IV  NOT_1258(g9529,I14672);
  IV  NOT_1259(g4164,I7311);
  IV  NOT_1260(g10538,I16181);
  IV  NOT_1261(g4233,g3698);
  IV  NOT_1262(g5424,I8865);
  IV  NOT_1263(g9348,I14549);
  IV  NOT_1264(I11326,g6660);
  IV  NOT_1265(I13949,g8451);
  IV  NOT_1266(g6403,g6128);
  IV  NOT_1267(I13326,g8203);
  IV  NOT_1268(I9804,g5417);
  IV  NOT_1269(g6145,I9860);
  IV  NOT_1270(g2859,I5995);
  IV  NOT_1271(g3997,I7131);
  IV  NOT_1272(I15510,g10035);
  IV  NOT_1273(g9355,I14570);
  IV  NOT_1274(I9792,g5403);
  IV  NOT_1275(I6832,g2909);
  IV  NOT_1276(g4454,g3914);
  IV  NOT_1277(g8033,I12875);
  IV  NOT_1278(g11510,I17549);
  IV  NOT_1279(g6191,g5446);
  IV  NOT_1280(g7569,I12029);
  IV  NOT_1281(g5672,I9177);
  IV  NOT_1282(g4296,I7559);
  IV  NOT_1283(I11904,g6902);
  IV  NOT_1284(I10633,g6015);
  IV  NOT_1285(I10898,g6735);
  IV  NOT_1286(g5231,g4640);
  IV  NOT_1287(I17318,g11340);
  IV  NOT_1288(g3332,I6513);
  IV  NOT_1289(I11252,g6542);
  IV  NOT_1290(g10241,g10192);
  IV  NOT_1291(g9260,g8892);
  IV  NOT_1292(g6695,I10666);
  IV  NOT_1293(I10719,g6003);
  IV  NOT_1294(I13621,g8315);
  IV  NOT_1295(g5643,I9090);
  IV  NOT_1296(g3353,g3121);
  IV  NOT_1297(I7735,g3759);
  IV  NOT_1298(I6507,g2808);
  IV  NOT_1299(I14191,g8795);
  IV  NOT_1300(g8096,I12953);
  IV  NOT_1301(g2248,g99);
  IV  NOT_1302(g11578,I17616);
  IV  NOT_1303(g2342,I5406);
  IV  NOT_1304(I7782,g3775);
  IV  NOT_1305(g6107,I9776);
  IV  NOT_1306(I17540,g11498);
  IV  NOT_1307(I12857,g7638);
  IV  NOT_1308(g11014,I16735);
  IV  NOT_1309(g6307,I10180);
  IV  NOT_1310(g3744,g3307);
  IV  NOT_1311(g6536,I10456);
  IV  NOT_1312(I4883,g581);
  IV  NOT_1313(g5205,g4366);
  IV  NOT_1314(I15586,g10159);
  IV  NOT_1315(I8880,g4537);
  IV  NOT_1316(g2255,I5276);
  IV  NOT_1317(I5728,g2084);
  IV  NOT_1318(g7688,g7148);
  IV  NOT_1319(I12793,g7619);
  IV  NOT_1320(g2481,g882);
  IV  NOT_1321(I9202,g4915);
  IV  NOT_1322(g8195,I13122);
  IV  NOT_1323(g7976,I12776);
  IV  NOT_1324(g8137,I13010);
  IV  NOT_1325(g8891,I14239);
  IV  NOT_1326(g8337,I13391);
  IV  NOT_1327(g10235,g10189);
  IV  NOT_1328(g4012,I7154);
  IV  NOT_1329(I11183,g6507);
  IV  NOT_1330(I16193,g10485);
  IV  NOT_1331(g11442,I17377);
  IV  NOT_1332(g2097,I4935);
  IV  NOT_1333(I12765,g7638);
  IV  NOT_1334(g10683,g10612);
  IV  NOT_1335(g5742,I9308);
  IV  NOT_1336(g2726,g2021);
  IV  NOT_1337(g4412,I7746);
  IV  NOT_1338(I11397,g6713);
  IV  NOT_1339(I13397,g8138);
  IV  NOT_1340(g2154,I5067);
  IV  NOT_1341(g6016,I9632);
  IV  NOT_1342(I12690,g7555);
  IV  NOT_1343(g4189,I7384);
  IV  NOT_1344(I5070,g1194);
  IV  NOT_1345(g2960,I6173);
  IV  NOT_1346(I10861,g6694);
  IV  NOT_1347(I10573,g5980);
  IV  NOT_1348(I9567,g5556);
  IV  NOT_1349(g8807,I14140);
  IV  NOT_1350(I14573,g9029);
  IV  NOT_1351(g4888,I8237);
  IV  NOT_1352(g7126,I11367);
  IV  NOT_1353(I13933,g8505);
  IV  NOT_1354(I17377,g11412);
  IV  NOT_1355(g7326,I11626);
  IV  NOT_1356(I10045,g5727);
  IV  NOT_1357(g6115,I9798);
  IV  NOT_1358(g6251,I10012);
  IV  NOT_1359(g4171,I7330);
  IV  NOT_1360(g6315,I10204);
  IV  NOT_1361(g6811,I10843);
  IV  NOT_1362(I15275,g9994);
  IV  NOT_1363(g4371,I7674);
  IV  NOT_1364(I14045,g8603);
  IV  NOT_1365(I17739,g11641);
  IV  NOT_1366(g4429,I7779);
  IV  NOT_1367(g4787,g3423);
  IV  NOT_1368(I8982,g4728);
  IV  NOT_1369(g11041,I16784);
  IV  NOT_1370(g10882,I16616);
  IV  NOT_1371(g5754,I9332);
  IV  NOT_1372(I9776,g5353);
  IV  NOT_1373(I10099,g5800);
  IV  NOT_1374(I16475,g10765);
  IV  NOT_1375(g6447,g6166);
  IV  NOT_1376(I10388,g5830);
  IV  NOT_1377(I8234,g4232);
  IV  NOT_1378(g7760,I12445);
  IV  NOT_1379(I14388,g8924);
  IV  NOT_1380(I8328,g4801);
  IV  NOT_1381(I17146,g11305);
  IV  NOT_1382(I16863,g10972);
  IV  NOT_1383(g3092,g2181);
  IV  NOT_1384(I14701,g9291);
  IV  NOT_1385(I10251,g6126);
  IV  NOT_1386(I14534,g9290);
  IV  NOT_1387(g4281,g3586);
  IV  NOT_1388(I9965,g5493);
  IV  NOT_1389(g5613,g4840);
  IV  NOT_1390(g6874,I10958);
  IV  NOT_1391(g8142,I13023);
  IV  NOT_1392(g2112,g639);
  IV  NOT_1393(g8342,I13406);
  IV  NOT_1394(g2218,g85);
  IV  NOT_1395(I15983,g10414);
  IV  NOT_1396(g2267,I5304);
  IV  NOT_1397(I17698,g11616);
  IV  NOT_1398(g11035,I16766);
  IV  NOT_1399(g8255,g7986);
  IV  NOT_1400(g8081,g8000);
  IV  NOT_1401(g8481,g8324);
  IV  NOT_1402(g2001,g814);
  IV  NOT_1403(g7608,I12174);
  IV  NOT_1404(g7924,g7470);
  IV  NOT_1405(I5406,g898);
  IV  NOT_1406(g7220,I11456);
  IV  NOT_1407(g5572,I8989);
  IV  NOT_1408(g5862,I9479);
  IV  NOT_1409(I12245,g7093);
  IV  NOT_1410(g7779,I12502);
  IV  NOT_1411(I4780,g872);
  IV  NOT_1412(I6040,g2216);
  IV  NOT_1413(g6595,I10563);
  IV  NOT_1414(g10584,g10522);
  IV  NOT_1415(I15517,g10051);
  IV  NOT_1416(I13574,g8360);
  IV  NOT_1417(g2329,I5383);
  IV  NOT_1418(g8354,I13442);
  IV  NOT_1419(I14140,g8717);
  IV  NOT_1420(g7023,I11166);
  IV  NOT_1421(I7952,g3664);
  IV  NOT_1422(g4963,I8337);
  IV  NOT_1423(g10206,g10178);
  IV  NOT_1424(I5801,g1984);
  IV  NOT_1425(I7276,g2861);
  IV  NOT_1426(g9670,I14799);
  IV  NOT_1427(I16781,g10893);
  IV  NOT_1428(g4791,I8161);
  IV  NOT_1429(g7977,I12779);
  IV  NOT_1430(g2828,I5940);
  IV  NOT_1431(g6272,I10075);
  IV  NOT_1432(I16236,g10535);
  IV  NOT_1433(g3262,I6432);
  IV  NOT_1434(g2727,g2022);
  IV  NOT_1435(g3736,I6924);
  IV  NOT_1436(g5534,g4545);
  IV  NOT_1437(g5729,I9279);
  IV  NOT_1438(g7361,I11731);
  IV  NOT_1439(g10114,I15350);
  IV  NOT_1440(I16175,g10488);
  IV  NOT_1441(g9813,I14948);
  IV  NOT_1442(I15193,g9968);
  IV  NOT_1443(g6417,g6136);
  IV  NOT_1444(I13051,g8060);
  IV  NOT_1445(I15362,g9987);
  IV  NOT_1446(g6935,I11065);
  IV  NOT_1447(g11193,g11112);
  IV  NOT_1448(g7051,I11232);
  IV  NOT_1449(g10107,I15341);
  IV  NOT_1450(I11756,g7191);
  IV  NOT_1451(g2221,I5198);
  IV  NOT_1452(g3076,I6282);
  IV  NOT_1453(I13592,g8362);
  IV  NOT_1454(g8783,g8746);
  IV  NOT_1455(I15523,g10058);
  IV  NOT_1456(g7327,I11629);
  IV  NOT_1457(I12232,g7072);
  IV  NOT_1458(I6528,g3274);
  IV  NOT_1459(I16264,g10557);
  IV  NOT_1460(g8979,I14358);
  IV  NOT_1461(I16790,g10900);
  IV  NOT_1462(I8490,g4526);
  IV  NOT_1463(g4201,I7420);
  IV  NOT_1464(I6648,g2635);
  IV  NOT_1465(g8218,g7826);
  IV  NOT_1466(I9658,g5150);
  IV  NOT_1467(g8312,I13320);
  IV  NOT_1468(I7546,g4105);
  IV  NOT_1469(g6128,I9829);
  IV  NOT_1470(g6629,I10584);
  IV  NOT_1471(g5885,g5361);
  IV  NOT_1472(g10345,I15801);
  IV  NOT_1473(g7999,I12825);
  IV  NOT_1474(g7146,I11391);
  IV  NOT_1475(g5660,I9141);
  IV  NOT_1476(I5445,g922);
  IV  NOT_1477(g6330,I10221);
  IV  NOT_1478(g7346,I11686);
  IV  NOT_1479(I10162,g5943);
  IV  NOT_1480(g7633,I12239);
  IV  NOT_1481(g4049,g3144);
  IV  NOT_1482(g3375,I6569);
  IV  NOT_1483(g8001,I12829);
  IV  NOT_1484(I12261,g7078);
  IV  NOT_1485(g4449,g4144);
  IV  NOT_1486(g3722,I6894);
  IV  NOT_1487(I8456,g4472);
  IV  NOT_1488(g7103,I11338);
  IV  NOT_1489(g5903,I9536);
  IV  NOT_1490(g4575,g3880);
  IV  NOT_1491(g10848,I16546);
  IV  NOT_1492(g11475,I17466);
  IV  NOT_1493(g8293,I13233);
  IV  NOT_1494(g8129,g8015);
  IV  NOT_1495(I6010,g2256);
  IV  NOT_1496(g2068,I4866);
  IV  NOT_1497(I11152,g6469);
  IV  NOT_1498(g8329,I13367);
  IV  NOT_1499(g10141,I15421);
  IV  NOT_1500(g7696,g7148);
  IV  NOT_1501(g10804,I16514);
  IV  NOT_1502(g6800,I10810);
  IV  NOT_1503(g4098,I7240);
  IV  NOT_1504(g3500,I6690);
  IV  NOT_1505(I15437,g10050);
  IV  NOT_1506(I16209,g10452);
  IV  NOT_1507(I8851,g4498);
  IV  NOT_1508(I11731,g7021);
  IV  NOT_1509(g8828,g8744);
  IV  NOT_1510(g11437,I17362);
  IV  NOT_1511(g2677,g2034);
  IV  NOT_1512(g10263,g10127);
  IV  NOT_1513(g7753,I12424);
  IV  NOT_1514(I9981,g5514);
  IV  NOT_1515(g8727,g8592);
  IV  NOT_1516(g5679,I9194);
  IV  NOT_1517(g7508,g6950);
  IV  NOT_1518(g3384,g3143);
  IV  NOT_1519(g10332,I15782);
  IV  NOT_1520(g6213,g5426);
  IV  NOT_1521(g8592,I13837);
  IV  NOT_1522(g7944,g7410);
  IV  NOT_1523(I15347,g9995);
  IV  NOT_1524(g7072,I11293);
  IV  NOT_1525(I15253,g9987);
  IV  NOT_1526(g10135,I15403);
  IV  NOT_1527(I12445,g7521);
  IV  NOT_1528(g11347,I17164);
  IV  NOT_1529(g4896,I8253);
  IV  NOT_1530(I7906,g3907);
  IV  NOT_1531(g2349,I5421);
  IV  NOT_1532(g7043,I11214);
  IV  NOT_1533(I12499,g7725);
  IV  NOT_1534(I11405,g6627);
  IV  NOT_1535(g5288,g4438);
  IV  NOT_1536(g9341,I14528);
  IV  NOT_1537(g3424,g2896);
  IV  NOT_1538(I9132,g4893);
  IV  NOT_1539(g10361,g10268);
  IV  NOT_1540(g3737,g2834);
  IV  NOT_1541(g7443,I11841);
  IV  NOT_1542(I9332,g4935);
  IV  NOT_1543(g9525,g9257);
  IV  NOT_1544(I9153,g5027);
  IV  NOT_1545(I9680,g5194);
  IV  NOT_1546(I10147,g5697);
  IV  NOT_1547(I6343,g1963);
  IV  NOT_1548(I10355,g6003);
  IV  NOT_1549(g7116,I11351);
  IV  NOT_1550(g5805,I9409);
  IV  NOT_1551(g5916,I9550);
  IV  NOT_1552(g7316,I11596);
  IV  NOT_1553(g2198,g668);
  IV  NOT_1554(I6282,g2231);
  IV  NOT_1555(g4268,I7523);
  IV  NOT_1556(I7771,g3418);
  IV  NOT_1557(I16607,g10787);
  IV  NOT_1558(g2855,I5989);
  IV  NOT_1559(g4362,I7651);
  IV  NOT_1560(I11929,g6901);
  IV  NOT_1561(I14355,g8948);
  IV  NOT_1562(I12989,g8043);
  IV  NOT_1563(g11351,I17170);
  IV  NOT_1564(g3077,g2213);
  IV  NOT_1565(g5422,g4470);
  IV  NOT_1566(g7034,I11191);
  IV  NOT_1567(I10825,g6588);
  IV  NOT_1568(g4419,I7763);
  IV  NOT_1569(I9744,g5263);
  IV  NOT_1570(I12056,g6929);
  IV  NOT_1571(I10370,g5857);
  IV  NOT_1572(g6166,I9893);
  IV  NOT_1573(g8624,g8486);
  IV  NOT_1574(g3523,g2971);
  IV  NOT_1575(I14370,g8954);
  IV  NOT_1576(g8953,I14312);
  IV  NOT_1577(I10858,g6688);
  IV  NOT_1578(I13020,g8049);
  IV  NOT_1579(I13583,g8344);
  IV  NOT_1580(g4452,g3365);
  IV  NOT_1581(I8872,g4529);
  IV  NOT_1582(I15063,g9699);
  IV  NOT_1583(g2241,g722);
  IV  NOT_1584(g7147,I11394);
  IV  NOT_1585(g6056,g5426);
  IV  NOT_1586(g5947,I9585);
  IV  NOT_1587(g7347,I11689);
  IV  NOT_1588(g11063,g10974);
  IV  NOT_1589(I11046,g6635);
  IV  NOT_1590(I10996,g6786);
  IV  NOT_1591(I12271,g7218);
  IV  NOT_1592(g7681,g7148);
  IV  NOT_1593(g6649,I10610);
  IV  NOT_1594(I8989,g4746);
  IV  NOT_1595(g8677,I13962);
  IV  NOT_1596(g110,I4786);
  IV  NOT_1597(I10367,g6234);
  IV  NOT_1598(I10394,g5824);
  IV  NOT_1599(I9901,g5557);
  IV  NOT_1600(g7697,g7101);
  IV  NOT_1601(I14367,g8953);
  IV  NOT_1602(I14394,g8884);
  IV  NOT_1603(I16641,g10864);
  IV  NOT_1604(g3742,I6929);
  IV  NOT_1605(g7914,g7651);
  IV  NOT_1606(g8576,I13819);
  IV  NOT_1607(g2524,g986);
  IV  NOT_1608(g7210,I11440);
  IV  NOT_1609(g4728,I8080);
  IV  NOT_1610(I16292,g10551);
  IV  NOT_1611(g2644,g1990);
  IV  NOT_1612(g6698,I10671);
  IV  NOT_1613(g4730,g3546);
  IV  NOT_1614(g8716,g8576);
  IV  NOT_1615(I17546,g11500);
  IV  NOT_1616(g8149,I13036);
  IV  NOT_1617(g10947,I16708);
  IV  NOT_1618(g4504,I7899);
  IV  NOT_1619(I11357,g6594);
  IV  NOT_1620(g6964,g6509);
  IV  NOT_1621(g8349,I13427);
  IV  NOT_1622(g2119,I5031);
  IV  NOT_1623(g5095,I8465);
  IV  NOT_1624(g6260,I10039);
  IV  NOT_1625(g5037,I8414);
  IV  NOT_1626(I13357,g8125);
  IV  NOT_1627(I12199,g7278);
  IV  NOT_1628(g4185,I7372);
  IV  NOT_1629(I7244,g3226);
  IV  NOT_1630(g9311,I14506);
  IV  NOT_1631(g11422,I17321);
  IV  NOT_1632(I11743,g7035);
  IV  NOT_1633(I13105,g7929);
  IV  NOT_1634(g5653,I9120);
  IV  NOT_1635(g4385,I7710);
  IV  NOT_1636(g7413,g7197);
  IV  NOT_1637(g5102,I8476);
  IV  NOT_1638(g2258,I5289);
  IV  NOT_1639(I14319,g8816);
  IV  NOT_1640(g2352,I5430);
  IV  NOT_1641(g2818,I5922);
  IV  NOT_1642(I7140,g2641);
  IV  NOT_1643(g6063,g5446);
  IV  NOT_1644(I12529,g7589);
  IV  NOT_1645(I5940,g2175);
  IV  NOT_1646(g2867,I6007);
  IV  NOT_1647(I16635,g10862);
  IV  NOT_1648(g10463,I15980);
  IV  NOT_1649(g11208,g11077);
  IV  NOT_1650(g4470,I7843);
  IV  NOT_1651(g8198,I13131);
  IV  NOT_1652(g4897,I8256);
  IV  NOT_1653(g8747,I14040);
  IV  NOT_1654(I7478,g3566);
  IV  NOT_1655(g5719,I9259);
  IV  NOT_1656(g4425,I7771);
  IV  NOT_1657(I12843,g7683);
  IV  NOT_1658(I15542,g10065);
  IV  NOT_1659(g10972,I16717);
  IV  NOT_1660(g10033,I15235);
  IV  NOT_1661(I5388,g889);
  IV  NOT_1662(g10234,g10188);
  IV  NOT_1663(I7435,g3459);
  IV  NOT_1664(g7936,g7712);
  IV  NOT_1665(g11542,g11519);
  IV  NOT_1666(g11453,I17416);
  IV  NOT_1667(g5752,I9326);
  IV  NOT_1668(I6094,g2110);
  IV  NOT_1669(I13803,g8476);
  IV  NOT_1670(g3044,I6256);
  IV  NOT_1671(g2211,g153);
  IV  NOT_1672(I14540,g9310);
  IV  NOT_1673(g6279,I10096);
  IV  NOT_1674(g2186,g90);
  IV  NOT_1675(g7317,I11599);
  IV  NOT_1676(g6720,I10713);
  IV  NOT_1677(I8253,g4637);
  IV  NOT_1678(g6118,I9807);
  IV  NOT_1679(g3983,g3222);
  IV  NOT_1680(g11614,I17662);
  IV  NOT_1681(g7601,I12153);
  IV  NOT_1682(I5430,g916);
  IV  NOT_1683(g5265,g4362);
  IV  NOT_1684(g11436,I17359);
  IV  NOT_1685(g3862,g2920);
  IV  NOT_1686(g5042,g4840);
  IV  NOT_1687(I15320,g10013);
  IV  NOT_1688(g9832,I14989);
  IV  NOT_1689(g6652,I10613);
  IV  NOT_1690(g4678,g3546);
  IV  NOT_1691(g6057,g5446);
  IV  NOT_1692(g6843,I10901);
  IV  NOT_1693(I15530,g10107);
  IV  NOT_1694(g11073,g10913);
  IV  NOT_1695(g4331,I7606);
  IV  NOT_1696(g3543,g3101);
  IV  NOT_1697(g2170,g30);
  IV  NOT_1698(g2614,g1994);
  IV  NOT_1699(g7775,I12490);
  IV  NOT_1700(g11593,I17633);
  IV  NOT_1701(g7922,I12712);
  IV  NOT_1702(g2125,I5053);
  IV  NOT_1703(g8319,I13341);
  IV  NOT_1704(g11346,I17161);
  IV  NOT_1705(I15565,g10101);
  IV  NOT_1706(g2821,I5929);
  IV  NOT_1707(g9507,g9268);
  IV  NOT_1708(I15464,g10094);
  IV  NOT_1709(I6965,g2880);
  IV  NOT_1710(I10120,g6248);
  IV  NOT_1711(g4766,g3440);
  IV  NOT_1712(I11662,g7033);
  IV  NOT_1713(I10739,g5942);
  IV  NOT_1714(g4087,I7220);
  IV  NOT_1715(g4105,I7249);
  IV  NOT_1716(g8152,I13043);
  IV  NOT_1717(g10421,g10331);
  IV  NOT_1718(I16537,g10721);
  IV  NOT_1719(g8352,I13436);
  IV  NOT_1720(g4305,g4013);
  IV  NOT_1721(g6971,g6517);
  IV  NOT_1722(I13027,g8051);
  IV  NOT_1723(I12258,g7103);
  IV  NOT_1724(g3729,I6907);
  IV  NOT_1725(I6264,g2118);
  IV  NOT_1726(I16108,g10383);
  IV  NOT_1727(g6686,I10651);
  IV  NOT_1728(g10163,I15485);
  IV  NOT_1729(g8717,I14010);
  IV  NOT_1730(g11034,I16763);
  IV  NOT_1731(g7460,g7148);
  IV  NOT_1732(g7597,I12133);
  IV  NOT_1733(g5296,g4444);
  IV  NOT_1734(I11249,g6541);
  IV  NOT_1735(I5638,g936);
  IV  NOT_1736(I14645,g9088);
  IV  NOT_1737(I16283,g10538);
  IV  NOT_1738(g2083,g139);
  IV  NOT_1739(I6360,g2261);
  IV  NOT_1740(g4748,g3546);
  IV  NOT_1741(I16492,g10773);
  IV  NOT_1742(I13482,g8193);
  IV  NOT_1743(I5308,g97);
  IV  NOT_1744(I11710,g7020);
  IV  NOT_1745(g7784,I12517);
  IV  NOT_1746(I4992,g1170);
  IV  NOT_1747(g4755,g3440);
  IV  NOT_1748(g10541,I16190);
  IV  NOT_1749(I10698,g5856);
  IV  NOT_1750(g6121,I9816);
  IV  NOT_1751(I15409,g10065);
  IV  NOT_1752(I7002,g2907);
  IV  NOT_1753(g8186,I13109);
  IV  NOT_1754(g10473,g10380);
  IV  NOT_1755(g4226,g3698);
  IV  NOT_1756(I11204,g6523);
  IV  NOT_1757(g6670,I10633);
  IV  NOT_1758(I7402,g4121);
  IV  NOT_1759(g11409,I17268);
  IV  NOT_1760(I6996,g2904);
  IV  NOT_1761(g3946,I7099);
  IV  NOT_1762(I13779,g8514);
  IV  NOT_1763(I7236,g3219);
  IV  NOT_1764(I15635,g10185);
  IV  NOT_1765(I16982,g11088);
  IV  NOT_1766(g8599,g8546);
  IV  NOT_1767(g7995,I12817);
  IV  NOT_1768(g2790,g2276);
  IV  NOT_1769(g11408,I17265);
  IV  NOT_1770(g7079,I11312);
  IV  NOT_1771(g11635,I17719);
  IV  NOT_1772(I11778,g7210);
  IV  NOT_1773(g3903,I7070);
  IV  NOT_1774(g5012,I8388);
  IV  NOT_1775(g9100,g8892);
  IV  NOT_1776(g8274,I13194);
  IV  NOT_1777(I10427,g5839);
  IV  NOT_1778(g7479,I11873);
  IV  NOT_1779(g8426,I13592);
  IV  NOT_1780(g1994,g794);
  IV  NOT_1781(g4445,I7803);
  IV  NOT_1782(g6253,I10018);
  IV  NOT_1783(g2061,g1828);
  IV  NOT_1784(g2187,g746);
  IV  NOT_1785(g6938,I11068);
  IV  NOT_1786(g4173,I7336);
  IV  NOT_1787(g6813,I10849);
  IV  NOT_1788(g4373,I7680);
  IV  NOT_1789(I11786,g7246);
  IV  NOT_1790(I16796,g11016);
  IV  NOT_1791(g10535,I16172);
  IV  NOT_1792(g4491,g3546);
  IV  NOT_1793(g8125,I12986);
  IV  NOT_1794(g7190,I11412);
  IV  NOT_1795(g8325,I13357);
  IV  NOT_1796(I11647,g6925);
  IV  NOT_1797(g7390,g6847);
  IV  NOT_1798(I12878,g7638);
  IV  NOT_1799(g5888,g5102);
  IV  NOT_1800(I13945,g8488);
  IV  NOT_1801(I12171,g6885);
  IV  NOT_1802(g10121,I15371);
  IV  NOT_1803(g8984,I14373);
  IV  NOT_1804(g3436,g3144);
  IV  NOT_1805(g4369,I7668);
  IV  NOT_1806(g8280,I13212);
  IV  NOT_1807(I7556,g4080);
  IV  NOT_1808(g4602,I8011);
  IV  NOT_1809(g7501,I11879);
  IV  NOT_1810(I17450,g11450);
  IV  NOT_1811(g3378,I6572);
  IV  NOT_1812(g5787,I9383);
  IV  NOT_1813(I9424,g4963);
  IV  NOT_1814(I9795,g5404);
  IV  NOT_1815(I17315,g11393);
  IV  NOT_1816(g10344,I15798);
  IV  NOT_1817(I9737,g5258);
  IV  NOT_1818(g2904,I6065);
  IV  NOT_1819(g2200,g92);
  IV  NOT_1820(g6552,g5733);
  IV  NOT_1821(g7356,I11716);
  IV  NOT_1822(g2046,g1845);
  IV  NOT_1823(I17707,g11619);
  IV  NOT_1824(g4920,I8293);
  IV  NOT_1825(I5827,g2271);
  IV  NOT_1826(g2446,g1400);
  IV  NOT_1827(g4459,I7820);
  IV  NOT_1828(I17202,g11322);
  IV  NOT_1829(g3335,I6520);
  IV  NOT_1830(I13233,g8265);
  IV  NOT_1831(g8483,g8332);
  IV  NOT_1832(g4767,I8123);
  IV  NOT_1833(I7064,g2984);
  IV  NOT_1834(g11575,g11561);
  IV  NOT_1835(g2003,g822);
  IV  NOT_1836(g5281,g4428);
  IV  NOT_1837(g3382,I6580);
  IV  NOT_1838(I9077,g4765);
  IV  NOT_1839(I7899,g3380);
  IV  NOT_1840(g4535,g3946);
  IV  NOT_1841(I8358,g4794);
  IV  NOT_1842(I6611,g2626);
  IV  NOT_1843(I8506,g4334);
  IV  NOT_1844(g2345,g1936);
  IV  NOT_1845(g10173,g10120);
  IV  NOT_1846(I17070,g11233);
  IV  NOT_1847(g8106,g7950);
  IV  NOT_1848(g11109,g10974);
  IV  NOT_1849(g8306,I13290);
  IV  NOT_1850(g2763,I5847);
  IV  NOT_1851(g2191,g1696);
  IV  NOT_1852(g2391,I5478);
  IV  NOT_1853(g6586,g5949);
  IV  NOT_1854(I12919,g8003);
  IV  NOT_1855(I6799,g2750);
  IV  NOT_1856(I11932,g6908);
  IV  NOT_1857(g3749,I6938);
  IV  NOT_1858(g8790,I14101);
  IV  NOT_1859(I9205,g5309);
  IV  NOT_1860(g11108,g10974);
  IV  NOT_1861(g2695,g2039);
  IV  NOT_1862(g9666,I14793);
  IV  NOT_1863(g8061,I12901);
  IV  NOT_1864(g5684,I9205);
  IV  NOT_1865(I8275,g4351);
  IV  NOT_1866(I8311,g4794);
  IV  NOT_1867(g4415,g3914);
  IV  NOT_1868(g5639,I9080);
  IV  NOT_1869(I14127,g8768);
  IV  NOT_1870(I17384,g11437);
  IV  NOT_1871(g7810,I12595);
  IV  NOT_1872(g7363,I11737);
  IV  NOT_1873(g10134,I15400);
  IV  NOT_1874(I7295,g3260);
  IV  NOT_1875(I11961,g7053);
  IV  NOT_1876(I16553,g10754);
  IV  NOT_1877(g5109,I8495);
  IV  NOT_1878(g5791,I9391);
  IV  NOT_1879(g3798,g3228);
  IV  NOT_1880(I13448,g8150);
  IV  NOT_1881(I9099,g5572);
  IV  NOT_1882(g2159,I5080);
  IV  NOT_1883(g7432,I11824);
  IV  NOT_1884(I14490,g8885);
  IV  NOT_1885(g6141,I9854);
  IV  NOT_1886(g8622,g8485);
  IV  NOT_1887(g6570,g5949);
  IV  NOT_1888(g6860,g6475);
  IV  NOT_1889(g7053,I11238);
  IV  NOT_1890(I11505,g6585);
  IV  NOT_1891(g9351,I14558);
  IV  NOT_1892(I5662,g563);
  IV  NOT_1893(g9875,I15036);
  IV  NOT_1894(g8427,I13595);
  IV  NOT_1895(I5067,g33);
  IV  NOT_1896(g9530,I14675);
  IV  NOT_1897(g6710,I10693);
  IV  NOT_1898(g5808,g5320);
  IV  NOT_1899(I5418,g907);
  IV  NOT_1900(g2858,I5992);
  IV  NOT_1901(I12598,g7628);
  IV  NOT_1902(I7194,g2629);
  IV  NOT_1903(I14376,g8959);
  IV  NOT_1904(I14385,g8890);
  IV  NOT_1905(g4203,I7426);
  IV  NOT_1906(I8985,g4733);
  IV  NOT_1907(I13717,g8354);
  IV  NOT_1908(g11381,I17206);
  IV  NOT_1909(g4721,g3546);
  IV  NOT_1910(g2016,g1361);
  IV  NOT_1911(I13212,g8195);
  IV  NOT_1912(g2757,I5837);
  IV  NOT_1913(g8446,I13636);
  IV  NOT_1914(g7568,I12026);
  IV  NOT_1915(g5759,I9341);
  IV  NOT_1916(I9754,g5271);
  IV  NOT_1917(I10888,g6333);
  IV  NOT_1918(g8514,I13711);
  IV  NOT_1919(I6802,g2751);
  IV  NOT_1920(g3632,I6799);
  IV  NOT_1921(g3095,g2482);
  IV  NOT_1922(g3037,g2135);
  IV  NOT_1923(g8003,I12835);
  IV  NOT_1924(I14888,g9454);
  IV  NOT_1925(I16252,g10515);
  IV  NOT_1926(g3437,I6654);
  IV  NOT_1927(I12817,g7692);
  IV  NOT_1928(I9273,g5091);
  IV  NOT_1929(I10671,g6045);
  IV  NOT_1930(I17695,g11614);
  IV  NOT_1931(g3102,g2482);
  IV  NOT_1932(I4924,g123);
  IV  NOT_1933(g3208,I6381);
  IV  NOT_1934(I12322,g7246);
  IV  NOT_1935(g7912,g7651);
  IV  NOT_1936(g8145,I13030);
  IV  NOT_1937(g8345,I13415);
  IV  NOT_1938(g2251,g731);
  IV  NOT_1939(g2642,g1988);
  IV  NOT_1940(I12159,g7243);
  IV  NOT_1941(g7357,I11719);
  IV  NOT_1942(g2047,g1857);
  IV  NOT_1943(I12532,g7594);
  IV  NOT_1944(I12901,g7984);
  IV  NOT_1945(g8191,I13114);
  IV  NOT_1946(g10927,g10827);
  IV  NOT_1947(g9884,I15063);
  IV  NOT_1948(g6158,I9883);
  IV  NOT_1949(g3719,g2920);
  IV  NOT_1950(I12783,g7590);
  IV  NOT_1951(g11390,I17219);
  IV  NOT_1952(I13723,g8359);
  IV  NOT_1953(g5865,I9486);
  IV  NOT_1954(g8695,I13978);
  IV  NOT_1955(I5847,g2275);
  IV  NOT_1956(I6901,g2818);
  IV  NOT_1957(I11149,g6468);
  IV  NOT_1958(g2874,I6022);
  IV  NOT_1959(g7929,g7519);
  IV  NOT_1960(g3752,I6947);
  IV  NOT_1961(I16673,g10782);
  IV  NOT_1962(I11433,g6424);
  IV  NOT_1963(I16847,g10886);
  IV  NOT_1964(I11387,g6672);
  IV  NOT_1965(g5604,I9032);
  IV  NOT_1966(I13433,g8181);
  IV  NOT_1967(g5098,g4840);
  IV  NOT_1968(g2654,g2012);
  IV  NOT_1969(I11620,g6840);
  IV  NOT_1970(g4188,I7381);
  IV  NOT_1971(g5498,I8919);
  IV  NOT_1972(I9712,g5230);
  IV  NOT_1973(g6587,g5827);
  IV  NOT_1974(g4388,I7719);
  IV  NOT_1975(g10491,I16108);
  IV  NOT_1976(g10903,g10809);
  IV  NOT_1977(I11097,g6748);
  IV  NOT_1978(I5421,g549);
  IV  NOT_1979(g8359,I13457);
  IV  NOT_1980(g6111,I9786);
  IV  NOT_1981(g6275,I10084);
  IV  NOT_1982(g6311,I10192);
  IV  NOT_1983(g4216,I7465);
  IV  NOT_1984(g10604,I16280);
  IV  NOT_1985(g9343,I14534);
  IV  NOT_1986(g8858,g8743);
  IV  NOT_1987(g4671,g3354);
  IV  NOT_1988(g2880,I6028);
  IV  NOT_1989(g4428,I7776);
  IV  NOT_1990(g2537,I5646);
  IV  NOT_1991(I10546,g5914);
  IV  NOT_1992(g5896,I9525);
  IV  NOT_1993(g4430,I7782);
  IV  NOT_1994(I14546,g9312);
  IV  NOT_1995(I7438,g3461);
  IV  NOT_1996(g3164,I6370);
  IV  NOT_1997(g3364,g3121);
  IV  NOT_1998(I7009,g2913);
  IV  NOT_1999(I10024,g5700);
  IV  NOT_2000(I8204,g3976);
  IV  NOT_2001(I12631,g7705);
  IV  NOT_2002(g8115,g7953);
  IV  NOT_2003(g4564,g3880);
  IV  NOT_2004(g8251,I13166);
  IV  NOT_2005(g8315,I13329);
  IV  NOT_2006(g2612,I5737);
  IV  NOT_2007(I15326,g10025);
  IV  NOT_2008(g2017,g1218);
  IV  NOT_2009(g6284,I10111);
  IV  NOT_2010(g2243,I5248);
  IV  NOT_2011(g8447,I13639);
  IV  NOT_2012(I6580,g3186);
  IV  NOT_2013(g3770,I6985);
  IV  NOT_2014(g6239,I9988);
  IV  NOT_2015(g10794,I16496);
  IV  NOT_2016(I15536,g10111);
  IV  NOT_2017(g10395,g10320);
  IV  NOT_2018(g5419,I8858);
  IV  NOT_2019(g9804,I14939);
  IV  NOT_2020(g10262,g10142);
  IV  NOT_2021(g7683,g7148);
  IV  NOT_2022(g11040,I16781);
  IV  NOT_2023(g10899,g10803);
  IV  NOT_2024(g6591,I10553);
  IV  NOT_2025(I11412,g6411);
  IV  NOT_2026(g5052,g4394);
  IV  NOT_2027(I13412,g8142);
  IV  NOT_2028(I5101,g1960);
  IV  NOT_2029(g8874,I14194);
  IV  NOT_2030(g3532,g3164);
  IV  NOT_2031(g7778,I12499);
  IV  NOT_2032(g2234,g87);
  IV  NOT_2033(g6853,I10917);
  IV  NOT_2034(I10126,g5682);
  IV  NOT_2035(I10659,g6038);
  IV  NOT_2036(I16574,g10821);
  IV  NOT_2037(g2629,g2001);
  IV  NOT_2038(g4638,g3354);
  IV  NOT_2039(g2328,g1882);
  IV  NOT_2040(I12289,g7142);
  IV  NOT_2041(I6968,g2881);
  IV  NOT_2042(g6420,I10334);
  IV  NOT_2043(g11621,I17681);
  IV  NOT_2044(g2130,I5057);
  IV  NOT_2045(g10191,I15551);
  IV  NOT_2046(g2542,g1868);
  IV  NOT_2047(I8973,g4488);
  IV  NOT_2048(g2330,g1891);
  IV  NOT_2049(g7735,I12384);
  IV  NOT_2050(I16311,g10584);
  IV  NOT_2051(g4308,g3863);
  IV  NOT_2052(I11228,g6471);
  IV  NOT_2053(I17231,g11303);
  IV  NOT_2054(g7782,I12511);
  IV  NOT_2055(g6559,g5758);
  IV  NOT_2056(I12571,g7509);
  IV  NOT_2057(g3012,I6247);
  IV  NOT_2058(I11011,g6340);
  IV  NOT_2059(I5751,g2296);
  IV  NOT_2060(g8595,I13840);
  IV  NOT_2061(g6931,I11055);
  IV  NOT_2062(g5728,I9276);
  IV  NOT_2063(g5486,g4395);
  IV  NOT_2064(I10296,g6242);
  IV  NOT_2065(I11716,g7026);
  IV  NOT_2066(g5730,I9282);
  IV  NOT_2067(g5504,g4419);
  IV  NOT_2068(g7949,g7422);
  IV  NOT_2069(g4217,I7468);
  IV  NOT_2070(g11183,I16950);
  IV  NOT_2071(I8123,g3630);
  IV  NOT_2072(g3990,g3121);
  IV  NOT_2073(g2554,I5672);
  IV  NOT_2074(g4758,g3586);
  IV  NOT_2075(g4066,I7191);
  IV  NOT_2076(g8272,I13188);
  IV  NOT_2077(I16592,g10781);
  IV  NOT_2078(g4589,I7996);
  IV  NOT_2079(g5185,g4682);
  IV  NOT_2080(g11397,I17234);
  IV  NOT_2081(g5881,g5361);
  IV  NOT_2082(g7627,I12223);
  IV  NOT_2083(g9094,g8892);
  IV  NOT_2084(I5041,g1179);
  IV  NOT_2085(I9135,g5198);
  IV  NOT_2086(g4466,I7833);
  IV  NOT_2087(g1992,g782);
  IV  NOT_2088(g6905,I11011);
  IV  NOT_2089(g8978,I14355);
  IV  NOT_2090(I5441,g919);
  IV  NOT_2091(g3371,g2837);
  IV  NOT_2092(g11062,g10937);
  IV  NOT_2093(I10060,g5752);
  IV  NOT_2094(g2213,g1110);
  IV  NOT_2095(g11509,I17546);
  IV  NOT_2096(g7998,I12822);
  IV  NOT_2097(g10247,I15639);
  IV  NOT_2098(g4165,g3164);
  IV  NOT_2099(g4365,g3880);
  IV  NOT_2100(I13627,g8326);
  IV  NOT_2101(g5425,g4300);
  IV  NOT_2102(g10389,g10307);
  IV  NOT_2103(g10926,g10827);
  IV  NOT_2104(I10855,g6685);
  IV  NOT_2105(I13959,g8451);
  IV  NOT_2106(I13379,g8133);
  IV  NOT_2107(g11508,I17543);
  IV  NOT_2108(g4711,I8061);
  IV  NOT_2109(g6100,I9759);
  IV  NOT_2110(I11112,g6445);
  IV  NOT_2111(g8982,I14367);
  IV  NOT_2112(g11634,I17716);
  IV  NOT_2113(g10612,I16286);
  IV  NOT_2114(g6300,I10159);
  IV  NOT_2115(g7603,I12159);
  IV  NOT_2116(g4055,g3144);
  IV  NOT_2117(g7039,I11204);
  IV  NOT_2118(I9749,g5266);
  IV  NOT_2119(g10388,g10305);
  IV  NOT_2120(I8351,g4794);
  IV  NOT_2121(g8234,g7826);
  IV  NOT_2122(g2902,I6061);
  IV  NOT_2123(g7439,I11833);
  IV  NOT_2124(g8128,I12993);
  IV  NOT_2125(g8328,I13364);
  IV  NOT_2126(g7850,I12647);
  IV  NOT_2127(g10534,I16169);
  IV  NOT_2128(g10098,I15332);
  IV  NOT_2129(I17456,g11453);
  IV  NOT_2130(g4333,g4144);
  IV  NOT_2131(I7837,g4158);
  IV  NOT_2132(g8330,I13370);
  IV  NOT_2133(g10251,g10195);
  IV  NOT_2134(g10272,g10168);
  IV  NOT_2135(g2090,I4920);
  IV  NOT_2136(g4774,I8136);
  IV  NOT_2137(I7462,g3721);
  IV  NOT_2138(I9798,g5415);
  IV  NOT_2139(I13096,g7925);
  IV  NOT_2140(g2166,I5101);
  IV  NOT_2141(g6750,I10759);
  IV  NOT_2142(g9264,I14477);
  IV  NOT_2143(I6424,g2462);
  IV  NOT_2144(g7702,g7079);
  IV  NOT_2145(g4196,I7405);
  IV  NOT_2146(g5678,I9191);
  IV  NOT_2147(I10503,g5858);
  IV  NOT_2148(I16413,g10663);
  IV  NOT_2149(g10462,I15977);
  IV  NOT_2150(g4396,I7735);
  IV  NOT_2151(g3138,I6356);
  IV  NOT_2152(g8800,I14123);
  IV  NOT_2153(I14503,g8920);
  IV  NOT_2154(I8410,g4283);
  IV  NOT_2155(g2056,I4859);
  IV  NOT_2156(I16691,g10788);
  IV  NOT_2157(g9360,I14579);
  IV  NOT_2158(g3109,g2482);
  IV  NOT_2159(g3791,I7014);
  IV  NOT_2160(g2456,g1397);
  IV  NOT_2161(g7919,g7512);
  IV  NOT_2162(g10032,I15232);
  IV  NOT_2163(g2529,I5638);
  IV  NOT_2164(g2649,g2005);
  IV  NOT_2165(g10140,I15418);
  IV  NOT_2166(g4780,g3440);
  IV  NOT_2167(I8839,g4484);
  IV  NOT_2168(g6040,I9655);
  IV  NOT_2169(g2348,I5418);
  IV  NOT_2170(I6077,g2349);
  IV  NOT_2171(g11574,g11561);
  IV  NOT_2172(g11452,I17413);
  IV  NOT_2173(g11047,I16802);
  IV  NOT_2174(g5682,I9199);
  IV  NOT_2175(g5766,I9346);
  IV  NOT_2176(g5105,I8487);
  IV  NOT_2177(g4509,I7906);
  IV  NOT_2178(g6440,g6150);
  IV  NOT_2179(g1976,g643);
  IV  NOT_2180(g11205,g11112);
  IV  NOT_2181(I6477,g2069);
  IV  NOT_2182(I9632,g5557);
  IV  NOT_2183(g7952,g7427);
  IV  NOT_2184(I15311,g10013);
  IV  NOT_2185(g9450,g9097);
  IV  NOT_2186(g5305,g4378);
  IV  NOT_2187(g5801,g5320);
  IV  NOT_2188(I5734,g2097);
  IV  NOT_2189(I6523,g2819);
  IV  NOT_2190(g2155,I5070);
  IV  NOT_2191(I4820,g865);
  IV  NOT_2192(I17243,g11396);
  IV  NOT_2193(g2355,I5435);
  IV  NOT_2194(g2851,I5979);
  IV  NOT_2195(I7249,g2833);
  IV  NOT_2196(I12559,g7477);
  IV  NOT_2197(I14315,g8815);
  IV  NOT_2198(I6643,g3008);
  IV  NOT_2199(g8213,g7826);
  IV  NOT_2200(I10819,g6706);
  IV  NOT_2201(g11311,I17100);
  IV  NOT_2202(I10910,g6703);
  IV  NOT_2203(I12424,g7635);
  IV  NOT_2204(I9102,g5586);
  IV  NOT_2205(I9208,g5047);
  IV  NOT_2206(g3707,g2920);
  IV  NOT_2207(I9302,g5576);
  IV  NOT_2208(I14910,g9532);
  IV  NOT_2209(g7616,I12196);
  IV  NOT_2210(g7561,I12015);
  IV  NOT_2211(g4067,I7194);
  IV  NOT_2212(g3759,I6958);
  IV  NOT_2213(I8278,g4495);
  IV  NOT_2214(I14257,g8805);
  IV  NOT_2215(g5748,I9320);
  IV  NOT_2216(I10979,g6565);
  IV  NOT_2217(g2964,I6193);
  IV  NOT_2218(g4418,I7760);
  IV  NOT_2219(I9869,g5405);
  IV  NOT_2220(g4467,g3829);
  IV  NOT_2221(I15072,g9713);
  IV  NOT_2222(I14979,g9671);
  IV  NOT_2223(g4290,g3586);
  IV  NOT_2224(I10111,g5754);
  IV  NOT_2225(I14055,g8650);
  IV  NOT_2226(g10871,I16583);
  IV  NOT_2227(g11051,I16814);
  IV  NOT_2228(I5992,g2195);
  IV  NOT_2229(g7004,I11143);
  IV  NOT_2230(I16583,g10848);
  IV  NOT_2231(g11072,g10913);
  IV  NOT_2232(I17773,g11650);
  IV  NOT_2233(I15592,g10163);
  IV  NOT_2234(I15756,g10266);
  IV  NOT_2235(g7527,g7148);
  IV  NOT_2236(I17268,g11351);
  IV  NOT_2237(I6742,g3326);
  IV  NOT_2238(I12544,g7669);
  IV  NOT_2239(g4093,g2965);
  IV  NOT_2240(I8282,g4770);
  IV  NOT_2241(g6151,I9872);
  IV  NOT_2242(g7764,I12457);
  IV  NOT_2243(g4256,g3664);
  IV  NOT_2244(g6648,I10607);
  IV  NOT_2245(g9777,g9474);
  IV  NOT_2246(g7546,I11970);
  IV  NOT_2247(I5080,g36);
  IV  NOT_2248(I15350,g10001);
  IV  NOT_2249(I10384,g5842);
  IV  NOT_2250(g10162,I15482);
  IV  NOT_2251(g3715,g2920);
  IV  NOT_2252(I9265,g5085);
  IV  NOT_2253(I16787,g10896);
  IV  NOT_2254(g11350,g11287);
  IV  NOT_2255(I5713,g2436);
  IV  NOT_2256(I15820,g10204);
  IV  NOT_2257(g5091,g4385);
  IV  NOT_2258(g8056,g7671);
  IV  NOT_2259(I13317,g8093);
  IV  NOT_2260(I12610,g7627);
  IV  NOT_2261(g4181,I7360);
  IV  NOT_2262(I6754,g2906);
  IV  NOT_2263(g8529,I13738);
  IV  NOT_2264(I14094,g8700);
  IV  NOT_2265(g4381,g3914);
  IV  NOT_2266(g7925,g7476);
  IV  NOT_2267(I9786,g5396);
  IV  NOT_2268(g2118,g1854);
  IV  NOT_2269(g8348,I13424);
  IV  NOT_2270(I12255,g7203);
  IV  NOT_2271(I6273,g2482);
  IV  NOT_2272(g2872,I6016);
  IV  NOT_2273(I16105,g10382);
  IV  NOT_2274(g10629,g10583);
  IV  NOT_2275(I10150,g5705);
  IV  NOT_2276(g5169,g4596);
  IV  NOT_2277(g4197,I7408);
  IV  NOT_2278(I10801,g6536);
  IV  NOT_2279(g8155,I13048);
  IV  NOT_2280(g11396,I17231);
  IV  NOT_2281(I13002,g8045);
  IV  NOT_2282(g8355,I13445);
  IV  NOT_2283(g10220,I15592);
  IV  NOT_2284(g5007,I8379);
  IV  NOT_2285(I13057,g7843);
  IV  NOT_2286(g2652,g2008);
  IV  NOT_2287(g2057,g754);
  IV  NOT_2288(g10628,I16307);
  IV  NOT_2289(I12678,g7376);
  IV  NOT_2290(I13128,g7976);
  IV  NOT_2291(g2843,I5963);
  IV  NOT_2292(g10911,I16685);
  IV  NOT_2293(g7320,I11608);
  IV  NOT_2294(g2989,g2135);
  IV  NOT_2295(g3539,g3015);
  IV  NOT_2296(g4263,g3586);
  IV  NOT_2297(I13245,g8269);
  IV  NOT_2298(I11626,g7042);
  IV  NOT_2299(I16769,g10894);
  IV  NOT_2300(g5718,I9256);
  IV  NOT_2301(I12460,g7569);
  IV  NOT_2302(I12939,g7977);
  IV  NOT_2303(g5767,I9349);
  IV  NOT_2304(I15691,g10233);
  IV  NOT_2305(I9296,g4908);
  IV  NOT_2306(I10018,g5862);
  IV  NOT_2307(I11299,g6727);
  IV  NOT_2308(I13323,g8203);
  IV  NOT_2309(I7176,g2623);
  IV  NOT_2310(I5976,g2186);
  IV  NOT_2311(g2549,g1386);
  IV  NOT_2312(I6572,g2853);
  IV  NOT_2313(I10526,g6161);
  IV  NOT_2314(g8063,I12907);
  IV  NOT_2315(g2834,I5952);
  IV  NOT_2316(g2971,g2046);
  IV  NOT_2317(g6172,I9901);
  IV  NOT_2318(g6278,I10093);
  IV  NOT_2319(g7617,I12199);
  IV  NOT_2320(I7405,g3861);
  IV  NOT_2321(g7906,I12694);
  IV  NOT_2322(g7789,I12532);
  IV  NOT_2323(g11405,I17258);
  IV  NOT_2324(g5261,g4640);
  IV  NOT_2325(g10591,I16258);
  IV  NOT_2326(I6543,g3186);
  IV  NOT_2327(g3362,I6546);
  IV  NOT_2328(g3419,g3104);
  IV  NOT_2329(I7829,g3425);
  IV  NOT_2330(g6667,I10630);
  IV  NOT_2331(g7516,g7148);
  IV  NOT_2332(g4562,I7973);
  IV  NOT_2333(g6343,I10248);
  IV  NOT_2334(g10754,I16439);
  IV  NOT_2335(g9353,I14564);
  IV  NOT_2336(g3052,I6264);
  IV  NOT_2337(g10355,I15829);
  IV  NOT_2338(g5415,I8848);
  IV  NOT_2339(g6282,I10105);
  IV  NOT_2340(g7771,I12478);
  IV  NOT_2341(g6566,g5791);
  IV  NOT_2342(I11737,g7027);
  IV  NOT_2343(g8279,I13209);
  IV  NOT_2344(g2121,I5041);
  IV  NOT_2345(g4631,g3820);
  IV  NOT_2346(I12875,g7638);
  IV  NOT_2347(g10825,I16537);
  IV  NOT_2348(I10917,g6732);
  IV  NOT_2349(I15583,g10157);
  IV  NOT_2350(g9802,g9490);
  IV  NOT_2351(g1999,g806);
  IV  NOT_2352(I11232,g6537);
  IV  NOT_2353(g4257,g3664);
  IV  NOT_2354(g6134,I9839);
  IV  NOT_2355(g5664,I9153);
  IV  NOT_2356(g8318,I13338);
  IV  NOT_2357(g8872,I14188);
  IV  NOT_2358(I9706,g5221);
  IV  NOT_2359(g2232,I5221);
  IV  NOT_2360(g10172,I15510);
  IV  NOT_2361(g11046,I16799);
  IV  NOT_2362(g3086,g2276);
  IV  NOT_2363(g5203,g4640);
  IV  NOT_2364(g2253,g100);
  IV  NOT_2365(g3728,I6904);
  IV  NOT_2366(g2813,I5913);
  IV  NOT_2367(I9029,g4781);
  IV  NOT_2368(g8989,I14388);
  IV  NOT_2369(I14077,g8758);
  IV  NOT_2370(I9171,g4902);
  IV  NOT_2371(g6555,g5740);
  IV  NOT_2372(I10706,g6080);
  IV  NOT_2373(I9371,g5075);
  IV  NOT_2374(g6804,I10822);
  IV  NOT_2375(I15787,g10269);
  IV  NOT_2376(I6414,g2342);
  IV  NOT_2377(g3730,g3015);
  IV  NOT_2378(g2909,I6080);
  IV  NOT_2379(I9956,g5485);
  IV  NOT_2380(I10689,g6059);
  IV  NOT_2381(g3385,g3121);
  IV  NOT_2382(I5383,g886);
  IV  NOT_2383(I15302,g10007);
  IV  NOT_2384(g11357,I17182);
  IV  NOT_2385(g7991,I12809);
  IV  NOT_2386(I6513,g2812);
  IV  NOT_2387(g2606,I5719);
  IV  NOT_2388(g10319,g10270);
  IV  NOT_2389(g4441,g3914);
  IV  NOT_2390(g6113,I9792);
  IV  NOT_2391(g6313,I10198);
  IV  NOT_2392(g7078,I11309);
  IV  NOT_2393(g7340,I11668);
  IV  NOT_2394(I10102,g5730);
  IV  NOT_2395(I16778,g10891);
  IV  NOT_2396(I13831,g8560);
  IV  NOT_2397(g10318,I15752);
  IV  NOT_2398(I8050,g4089);
  IV  NOT_2399(I13445,g8149);
  IV  NOT_2400(I5588,g1203);
  IV  NOT_2401(g8121,I12978);
  IV  NOT_2402(g10227,I15601);
  IV  NOT_2403(g7907,g7664);
  IV  NOT_2404(I6436,g2351);
  IV  NOT_2405(I6679,g2902);
  IV  NOT_2406(g8321,I13347);
  IV  NOT_2407(g4673,g4013);
  IV  NOT_2408(g6202,g5426);
  IV  NOT_2409(g8670,g8551);
  IV  NOT_2410(g5689,I9216);
  IV  NOT_2411(I8996,g4757);
  IV  NOT_2412(I9684,g5426);
  IV  NOT_2413(g7035,I11194);
  IV  NOT_2414(I15768,g10249);
  IV  NOT_2415(I9138,g5210);
  IV  NOT_2416(I9639,g5126);
  IV  NOT_2417(g7959,I12751);
  IV  NOT_2418(I10066,g5778);
  IV  NOT_2419(I9338,g5576);
  IV  NOT_2420(I10231,g6111);
  IV  NOT_2421(g8625,g8487);
  IV  NOT_2422(g7082,I11315);
  IV  NOT_2423(g2586,g1972);
  IV  NOT_2424(g5216,g4445);
  IV  NOT_2425(g10540,I16187);
  IV  NOT_2426(I17410,g11419);
  IV  NOT_2427(g6094,I9749);
  IV  NOT_2428(I11498,g6578);
  IV  NOT_2429(I12595,g7706);
  IV  NOT_2430(I16647,g10866);
  IV  NOT_2431(g10058,I15281);
  IV  NOT_2432(I16356,g10597);
  IV  NOT_2433(g4669,g4013);
  IV  NOT_2434(I8724,g4791);
  IV  NOT_2435(g6567,I10495);
  IV  NOT_2436(g5671,I9174);
  IV  NOT_2437(g4368,I7665);
  IV  NOT_2438(I11989,g6919);
  IV  NOT_2439(I17666,g11603);
  IV  NOT_2440(I10885,g6332);
  IV  NOT_2441(I8379,g4231);
  IV  NOT_2442(g3331,I6510);
  IV  NOT_2443(g10203,g10177);
  IV  NOT_2444(I14876,g9526);
  IV  NOT_2445(I11611,g6913);
  IV  NOT_2446(g7656,I12265);
  IV  NOT_2447(g4772,g3440);
  IV  NOT_2448(g3406,I6611);
  IV  NOT_2449(I11722,g7034);
  IV  NOT_2450(I7399,g4113);
  IV  NOT_2451(g10044,I15263);
  IV  NOT_2452(g3635,I6812);
  IV  NOT_2453(I6022,g2258);
  IV  NOT_2454(g4458,I7817);
  IV  NOT_2455(g2570,g207);
  IV  NOT_2456(g2860,I5998);
  IV  NOT_2457(g2341,I5403);
  IV  NOT_2458(g9262,I14473);
  IV  NOT_2459(g3682,g2920);
  IV  NOT_2460(g6593,I10557);
  IV  NOT_2461(I9759,g5344);
  IV  NOT_2462(g8519,I13726);
  IV  NOT_2463(g3105,g2482);
  IV  NOT_2464(g7915,g7473);
  IV  NOT_2465(g3305,I6474);
  IV  NOT_2466(g10281,g10162);
  IV  NOT_2467(g98,I4783);
  IV  NOT_2468(g2645,g1991);
  IV  NOT_2469(I8835,g4791);
  IV  NOT_2470(g5826,I9440);
  IV  NOT_2471(I12418,g7568);
  IV  NOT_2472(I12822,g7677);
  IV  NOT_2473(g10902,I16660);
  IV  NOT_2474(g10377,I15855);
  IV  NOT_2475(g8606,g8481);
  IV  NOT_2476(g7214,I11450);
  IV  NOT_2477(I6947,g2860);
  IV  NOT_2478(g10120,I15368);
  IV  NOT_2479(g4011,I7151);
  IV  NOT_2480(g9076,g8892);
  IV  NOT_2481(g5741,I9305);
  IV  NOT_2482(g3748,g2971);
  IV  NOT_2483(g4411,I7743);
  IV  NOT_2484(g4734,g3586);
  IV  NOT_2485(I11342,g6686);
  IV  NOT_2486(g9889,I15072);
  IV  NOT_2487(g7110,I11345);
  IV  NOT_2488(g6264,I10051);
  IV  NOT_2489(g7310,I11578);
  IV  NOT_2490(I6560,g2845);
  IV  NOT_2491(I7291,g3212);
  IV  NOT_2492(I8611,g4562);
  IV  NOT_2493(I10456,g5844);
  IV  NOT_2494(I15482,g10115);
  IV  NOT_2495(g5638,I9077);
  IV  NOT_2496(g3226,I6403);
  IV  NOT_2497(g6933,I11061);
  IV  NOT_2498(g7663,I12282);
  IV  NOT_2499(I11650,g6938);
  IV  NOT_2500(g10699,I16376);
  IV  NOT_2501(g2607,I5722);
  IV  NOT_2502(I12853,g7638);
  IV  NOT_2503(I16897,g10947);
  IV  NOT_2504(I5240,g64);
  IV  NOT_2505(g2962,I6183);
  IV  NOT_2506(g6521,I10437);
  IV  NOT_2507(I17084,g11249);
  IV  NOT_2508(g4474,g3820);
  IV  NOT_2509(g10290,I15694);
  IV  NOT_2510(g2158,I5077);
  IV  NOT_2511(g6050,I9677);
  IV  NOT_2512(g6641,I10598);
  IV  NOT_2513(I11198,g6521);
  IV  NOT_2514(I9498,g5081);
  IV  NOT_2515(I12589,g7571);
  IV  NOT_2516(g10698,I16373);
  IV  NOT_2517(g2506,g636);
  IV  NOT_2518(g6450,I10378);
  IV  NOT_2519(I6037,g2560);
  IV  NOT_2520(I17321,g11348);
  IV  NOT_2521(g5883,g5309);
  IV  NOT_2522(I10314,g6251);
  IV  NOT_2523(g7402,g6860);
  IV  NOT_2524(I6495,g2076);
  IV  NOT_2525(I9833,g5197);
  IV  NOT_2526(I17179,g11307);
  IV  NOT_2527(I11528,g6796);
  IV  NOT_2528(I6102,g2240);
  IV  NOT_2529(I16717,g10779);
  IV  NOT_2530(I17531,g11488);
  IV  NOT_2531(I7694,g3742);
  IV  NOT_2532(I11330,g6571);
  IV  NOT_2533(I6302,g2243);
  IV  NOT_2534(g3373,I6565);
  IV  NOT_2535(I15778,g10255);
  IV  NOT_2536(g7762,I12451);
  IV  NOT_2537(g3491,g2669);
  IV  NOT_2538(g4080,g2903);
  IV  NOT_2539(I5116,g40);
  IV  NOT_2540(g11081,I16856);
  IV  NOT_2541(I7852,g3438);
  IV  NOT_2542(I7923,g3394);
  IV  NOT_2543(g5758,I9338);
  IV  NOT_2544(g8141,I13020);
  IV  NOT_2545(g8570,I13803);
  IV  NOT_2546(g5066,I8436);
  IV  NOT_2547(g5589,I9001);
  IV  NOT_2548(g6724,I10719);
  IV  NOT_2549(g8341,I13403);
  IV  NOT_2550(I10054,g5728);
  IV  NOT_2551(g2275,g757);
  IV  NOT_2552(I9539,g5354);
  IV  NOT_2553(I9896,g5295);
  IV  NOT_2554(g4713,g3546);
  IV  NOT_2555(I10243,g5918);
  IV  NOT_2556(I11132,g6451);
  IV  NOT_2557(I11869,g6894);
  IV  NOT_2558(g7877,g7479);
  IV  NOT_2559(I7701,g3513);
  IV  NOT_2560(g3369,I6557);
  IV  NOT_2561(I5565,g1713);
  IV  NOT_2562(g3007,I6240);
  IV  NOT_2563(g9339,I14522);
  IV  NOT_2564(I15356,g10013);
  IV  NOT_2565(g7657,I12268);
  IV  NOT_2566(g6878,I10966);
  IV  NOT_2567(I15826,g10205);
  IV  NOT_2568(I6917,g2832);
  IV  NOT_2569(I15380,g10098);
  IV  NOT_2570(I4894,g258);
  IV  NOT_2571(g2174,g31);
  IV  NOT_2572(g3459,I6661);
  IV  NOT_2573(g6289,I10126);
  IV  NOT_2574(g9024,I14409);
  IV  NOT_2575(g2374,g591);
  IV  NOT_2576(I12616,g7534);
  IV  NOT_2577(I9162,g5035);
  IV  NOT_2578(g7556,I11992);
  IV  NOT_2579(I9268,g5305);
  IV  NOT_2580(I16723,g10851);
  IV  NOT_2581(g3767,I6976);
  IV  NOT_2582(g10547,I16206);
  IV  NOT_2583(g9424,g9076);
  IV  NOT_2584(g10895,I16647);
  IV  NOT_2585(I7886,g4076);
  IV  NOT_2586(I9362,g5013);
  IV  NOT_2587(g6835,I10885);
  IV  NOT_2588(g2985,I6217);
  IV  NOT_2589(g9809,I14944);
  IV  NOT_2590(g5827,I9443);
  IV  NOT_2591(g6882,I10974);
  IV  NOT_2592(g7928,g7508);
  IV  NOT_2593(I10156,g6100);
  IV  NOT_2594(I10655,g6036);
  IV  NOT_2595(I15672,g10132);
  IV  NOT_2596(g3582,g3164);
  IV  NOT_2597(I16387,g10629);
  IV  NOT_2598(I17334,g11360);
  IV  NOT_2599(g6271,I10072);
  IV  NOT_2600(I11225,g6534);
  IV  NOT_2601(g10226,I15598);
  IV  NOT_2602(I9452,g5085);
  IV  NOT_2603(g11182,I16947);
  IV  NOT_2604(g11651,I17755);
  IV  NOT_2605(g7064,I11269);
  IV  NOT_2606(I5210,g58);
  IV  NOT_2607(g2239,I5240);
  IV  NOT_2608(I10180,g6107);
  IV  NOT_2609(g9672,I14805);
  IV  NOT_2610(I13708,g8337);
  IV  NOT_2611(g5774,I9362);
  IV  NOT_2612(g7899,I12683);
  IV  NOT_2613(g3793,g2593);
  IV  NOT_2614(g7464,I11858);
  IV  NOT_2615(I12053,g6928);
  IV  NOT_2616(g8358,I13454);
  IV  NOT_2617(I12809,g7686);
  IV  NOT_2618(g7785,I12520);
  IV  NOT_2619(I16811,g10908);
  IV  NOT_2620(g10551,I16214);
  IV  NOT_2621(I6233,g2299);
  IV  NOT_2622(g2832,I5946);
  IV  NOT_2623(I12466,g7585);
  IV  NOT_2624(g3415,g3121);
  IV  NOT_2625(g3227,I6406);
  IV  NOT_2626(I7825,g3414);
  IV  NOT_2627(g6799,I10807);
  IV  NOT_2628(g2853,g2171);
  IV  NOT_2629(I11043,g6412);
  IV  NOT_2630(I6454,g2368);
  IV  NOT_2631(I13043,g8055);
  IV  NOT_2632(I17216,g11291);
  IV  NOT_2633(g2420,g237);
  IV  NOT_2634(g6674,I10639);
  IV  NOT_2635(I9486,g5066);
  IV  NOT_2636(g11513,I17558);
  IV  NOT_2637(I12177,g7259);
  IV  NOT_2638(g10127,I15383);
  IV  NOT_2639(g3664,g3209);
  IV  NOT_2640(g8275,I13197);
  IV  NOT_2641(g2507,I5584);
  IV  NOT_2642(g8311,I13317);
  IV  NOT_2643(g3246,g2482);
  IV  NOT_2644(I15448,g10056);
  IV  NOT_2645(g5509,g4739);
  IV  NOT_2646(g4326,g3863);
  IV  NOT_2647(I14694,g9259);
  IV  NOT_2648(I7408,g4125);
  IV  NOT_2649(g7237,I11477);
  IV  NOT_2650(g10490,I16105);
  IV  NOT_2651(I9185,g4915);
  IV  NOT_2652(I7336,g3997);
  IV  NOT_2653(g3721,I6891);
  IV  NOT_2654(g11505,I17534);
  IV  NOT_2655(I11602,g6833);
  IV  NOT_2656(I11810,g7246);
  IV  NOT_2657(g11404,I17255);
  IV  NOT_2658(g6132,I9833);
  IV  NOT_2659(g5662,I9147);
  IV  NOT_2660(I6553,g3186);
  IV  NOT_2661(I4850,g1958);
  IV  NOT_2662(g7844,I12631);
  IV  NOT_2663(I17543,g11499);
  IV  NOT_2664(I11068,g6426);
  IV  NOT_2665(I13068,g7906);
  IV  NOT_2666(g6680,I10643);
  IV  NOT_2667(g6209,I9956);
  IV  NOT_2668(g8985,I14376);
  IV  NOT_2669(I11879,g6893);
  IV  NOT_2670(g5994,I9612);
  IV  NOT_2671(g10889,I16629);
  IV  NOT_2672(I16850,g10905);
  IV  NOT_2673(I11970,g6918);
  IV  NOT_2674(g7394,I11778);
  IV  NOT_2675(I10557,g6197);
  IV  NOT_2676(g10354,I15826);
  IV  NOT_2677(g2905,I6068);
  IV  NOT_2678(g7089,I11322);
  IV  NOT_2679(g7731,I12376);
  IV  NOT_2680(g10888,I16626);
  IV  NOT_2681(g6802,I10816);
  IV  NOT_2682(g8239,g7826);
  IV  NOT_2683(g4183,I7366);
  IV  NOT_2684(g9273,I14490);
  IV  NOT_2685(g4608,g3829);
  IV  NOT_2686(g5816,I9424);
  IV  NOT_2687(I5922,g2170);
  IV  NOT_2688(I7465,g3726);
  IV  NOT_2689(g7966,I12762);
  IV  NOT_2690(g2100,I4948);
  IV  NOT_2691(I10278,g5815);
  IV  NOT_2692(g3940,g2920);
  IV  NOT_2693(g6558,I10484);
  IV  NOT_2694(I12009,g6915);
  IV  NOT_2695(I6888,g2960);
  IV  NOT_2696(I8262,g4636);
  IV  NOT_2697(I11967,g6911);
  IV  NOT_2698(g8020,I12862);
  IV  NOT_2699(I10286,g6237);
  IV  NOT_2700(g8420,I13574);
  IV  NOT_2701(I5060,g1191);
  IV  NOT_2702(g10931,g10827);
  IV  NOT_2703(g3388,I6590);
  IV  NOT_2704(I10039,g5718);
  IV  NOT_2705(I14306,g8812);
  IV  NOT_2706(I11459,g6488);
  IV  NOT_2707(g11433,I17350);
  IV  NOT_2708(g9572,I14709);
  IV  NOT_2709(g5685,I9208);
  IV  NOT_2710(g5197,I8611);
  IV  NOT_2711(g5700,I9237);
  IV  NOT_2712(g8794,I14109);
  IV  NOT_2713(g5397,I8835);
  IV  NOT_2714(g2750,I5818);
  IV  NOT_2715(I8889,g4553);
  IV  NOT_2716(g11620,I17678);
  IV  NOT_2717(g10190,I15548);
  IV  NOT_2718(I8476,g4577);
  IV  NOT_2719(g4361,I7648);
  IV  NOT_2720(I9766,g5348);
  IV  NOT_2721(I15811,g10200);
  IV  NOT_2722(g3428,I6639);
  IV  NOT_2723(I7096,g3186);
  IV  NOT_2724(I12454,g7544);
  IV  NOT_2725(I9087,g5113);
  IV  NOT_2726(I9105,g5589);
  IV  NOT_2727(I9305,g4970);
  IV  NOT_2728(I9801,g5416);
  IV  NOT_2729(g3430,I6643);
  IV  NOT_2730(g7814,I12607);
  IV  NOT_2731(I12712,g7441);
  IV  NOT_2732(g11646,I17742);
  IV  NOT_2733(g4051,I7166);
  IV  NOT_2734(I10601,g5996);
  IV  NOT_2735(I13010,g8047);
  IV  NOT_2736(g11343,I17152);
  IV  NOT_2737(I13918,g8451);
  IV  NOT_2738(I16379,g10598);
  IV  NOT_2739(g4127,I7276);
  IV  NOT_2740(g4451,g3638);
  IV  NOT_2741(I15971,g10408);
  IV  NOT_2742(g4327,I7600);
  IV  NOT_2743(I17265,g11352);
  IV  NOT_2744(g7350,I11698);
  IV  NOT_2745(g2040,g1786);
  IV  NOT_2746(g6574,I10514);
  IV  NOT_2747(I12907,g7959);
  IV  NOT_2748(I5995,g2196);
  IV  NOT_2749(I11079,g6649);
  IV  NOT_2750(g10546,I16203);
  IV  NOT_2751(g7038,I11201);
  IV  NOT_2752(I11444,g6653);
  IV  NOT_2753(I17416,g11420);
  IV  NOT_2754(g10211,I15583);
  IV  NOT_2755(g9534,I14687);
  IV  NOT_2756(g9961,I15162);
  IV  NOT_2757(g6714,g5867);
  IV  NOT_2758(g7438,g7232);
  IV  NOT_2759(g7773,I12484);
  IV  NOT_2760(I11599,g6832);
  IV  NOT_2761(g7009,I11152);
  IV  NOT_2762(g11369,I17194);
  IV  NOT_2763(g2123,I5047);
  IV  NOT_2764(I6639,g2632);
  IV  NOT_2765(g4346,I7625);
  IV  NOT_2766(g8515,I13714);
  IV  NOT_2767(g10088,I15317);
  IV  NOT_2768(I8285,g4771);
  IV  NOT_2769(I10937,g6552);
  IV  NOT_2770(I12239,g7073);
  IV  NOT_2771(I5840,g2432);
  IV  NOT_2772(I15368,g9990);
  IV  NOT_2773(I17510,g11481);
  IV  NOT_2774(I16742,g10857);
  IV  NOT_2775(g8100,g7947);
  IV  NOT_2776(I16944,g11079);
  IV  NOT_2777(g3910,g3015);
  IV  NOT_2778(I13086,g7924);
  IV  NOT_2779(g7769,I12472);
  IV  NOT_2780(I15412,g10075);
  IV  NOT_2781(g3638,I6821);
  IV  NOT_2782(I8139,g3681);
  IV  NOT_2783(g7212,I11444);
  IV  NOT_2784(g5723,I9265);
  IV  NOT_2785(I14884,g9454);
  IV  NOT_2786(g11412,I17277);
  IV  NOT_2787(I11817,g7246);
  IV  NOT_2788(I10168,g5982);
  IV  NOT_2789(g5101,I8473);
  IV  NOT_2790(g5817,I9427);
  IV  NOT_2791(I11322,g6652);
  IV  NOT_2792(g7918,g7505);
  IV  NOT_2793(g5301,g4373);
  IV  NOT_2794(g7967,I12765);
  IV  NOT_2795(g6262,I10045);
  IV  NOT_2796(I15229,g9968);
  IV  NOT_2797(g2351,I5427);
  IV  NOT_2798(I11159,g6478);
  IV  NOT_2799(g10700,I16379);
  IV  NOT_2800(g2648,I5765);
  IV  NOT_2801(I9491,g5072);
  IV  NOT_2802(g10126,I15380);
  IV  NOT_2803(I8024,g4117);
  IV  NOT_2804(I11901,g6897);
  IV  NOT_2805(I16802,g10902);
  IV  NOT_2806(g2530,I5641);
  IV  NOT_2807(g6736,I10739);
  IV  NOT_2808(I13125,g7975);
  IV  NOT_2809(g8750,I14045);
  IV  NOT_2810(I10666,g6042);
  IV  NOT_2811(g4508,g3946);
  IV  NOT_2812(g10250,g10136);
  IV  NOT_2813(g2655,g2013);
  IV  NOT_2814(g4944,g4430);
  IV  NOT_2815(g4240,g3664);
  IV  NOT_2816(I11783,g7246);
  IV  NOT_2817(I16793,g11014);
  IV  NOT_2818(I7342,g4011);
  IV  NOT_2819(I9602,g5013);
  IV  NOT_2820(g4472,I7847);
  IV  NOT_2821(I10015,g5641);
  IV  NOT_2822(I5704,g2056);
  IV  NOT_2823(g7993,I12813);
  IV  NOT_2824(I7255,g3227);
  IV  NOT_2825(g6076,I9717);
  IV  NOT_2826(I4906,g119);
  IV  NOT_2827(I11656,g7122);
  IV  NOT_2828(I6049,g2219);
  IV  NOT_2829(g5751,I9323);
  IV  NOT_2830(g3758,I6955);
  IV  NOT_2831(g3066,g2135);
  IV  NOT_2832(I8231,g4170);
  IV  NOT_2833(g4443,g3359);
  IV  NOT_2834(g10296,I15708);
  IV  NOT_2835(g8440,I13618);
  IV  NOT_2836(I11680,g7064);
  IV  NOT_2837(g8969,I14340);
  IV  NOT_2838(I17116,g11229);
  IV  NOT_2839(g2410,g1453);
  IV  NOT_2840(g9679,g9452);
  IV  NOT_2841(I7726,g3378);
  IV  NOT_2842(g6175,g5320);
  IV  NOT_2843(g4116,I7260);
  IV  NOT_2844(I7154,g2617);
  IV  NOT_2845(g8323,I13351);
  IV  NOT_2846(g6871,g6724);
  IV  NOT_2847(g2884,I6040);
  IV  NOT_2848(I7354,g4066);
  IV  NOT_2849(g2839,I5957);
  IV  NOT_2850(g3365,I6553);
  IV  NOT_2851(g3861,I7054);
  IV  NOT_2852(I6498,g2958);
  IV  NOT_2853(I17746,g11643);
  IV  NOT_2854(g3055,g2135);
  IV  NOT_2855(I5053,g1188);
  IV  NOT_2856(I15959,g10402);
  IV  NOT_2857(g6285,I10114);
  IV  NOT_2858(g11627,I17695);
  IV  NOT_2859(g7921,g7463);
  IV  NOT_2860(g10197,I15565);
  IV  NOT_2861(g5673,I9180);
  IV  NOT_2862(g4347,g3880);
  IV  NOT_2863(I8551,g4342);
  IV  NOT_2864(I10084,g5742);
  IV  NOT_2865(g2172,g43);
  IV  NOT_2866(g3333,g2779);
  IV  NOT_2867(I9415,g5047);
  IV  NOT_2868(g11112,I16897);
  IV  NOT_2869(I17237,g11394);
  IV  NOT_2870(g4681,g3546);
  IV  NOT_2871(g10870,I16580);
  IV  NOT_2872(g11050,I16811);
  IV  NOT_2873(I8499,g4330);
  IV  NOT_2874(I12577,g7532);
  IV  NOT_2875(g8151,g8036);
  IV  NOT_2876(g10527,g10462);
  IV  NOT_2877(g3774,I6999);
  IV  NOT_2878(g8351,I13433);
  IV  NOT_2879(I17340,g11366);
  IV  NOT_2880(g4533,I7938);
  IV  NOT_2881(I13017,g7848);
  IV  NOT_2882(I13364,g8221);
  IV  NOT_2883(I15386,g10101);
  IV  NOT_2884(g6184,I9915);
  IV  NOT_2885(g2235,g96);
  IV  NOT_2886(g2343,g1927);
  IV  NOT_2887(I12439,g7663);
  IV  NOT_2888(g5669,I9168);
  IV  NOT_2889(I10531,g6169);
  IV  NOT_2890(I17684,g11609);
  IV  NOT_2891(g6339,I10240);
  IV  NOT_2892(I14179,g8785);
  IV  NOT_2893(g4210,I7447);
  IV  NOT_2894(I14531,g9273);
  IV  NOT_2895(I7112,g3186);
  IV  NOT_2896(I17142,g11301);
  IV  NOT_2897(g11096,I16879);
  IV  NOT_2898(g7620,I12208);
  IV  NOT_2899(g4596,I8007);
  IV  NOT_2900(g3538,I6726);
  IV  NOT_2901(I6019,g2554);
  IV  NOT_2902(g4013,I7157);
  IV  NOT_2903(g6424,g6140);
  IV  NOT_2904(I16626,g10859);
  IV  NOT_2905(I10186,g6110);
  IV  NOT_2906(g6737,g6016);
  IV  NOT_2907(g10867,I16571);
  IV  NOT_2908(g2334,I5388);
  IV  NOT_2909(g10894,I16644);
  IV  NOT_2910(g6809,I10837);
  IV  NOT_2911(I10685,g6054);
  IV  NOT_2912(g5743,I9311);
  IV  NOT_2913(g4413,I7749);
  IV  NOT_2914(g5890,g5361);
  IV  NOT_2915(I11289,g6508);
  IV  NOT_2916(I6052,g2220);
  IV  NOT_2917(g2548,I5667);
  IV  NOT_2918(I14373,g8956);
  IV  NOT_2919(I11309,g6531);
  IV  NOT_2920(I5929,g2225);
  IV  NOT_2921(I13023,g8050);
  IV  NOT_2922(g8884,I14224);
  IV  NOT_2923(I16298,g10553);
  IV  NOT_2924(I13224,g8261);
  IV  NOT_2925(g7788,I12529);
  IV  NOT_2926(g6077,I9720);
  IV  NOT_2927(g11429,I17340);
  IV  NOT_2928(g5011,I8385);
  IV  NOT_2929(I16775,g10889);
  IV  NOT_2930(g3067,I6273);
  IV  NOT_2931(I13571,g8355);
  IV  NOT_2932(g10315,g10243);
  IV  NOT_2933(g5856,g5245);
  IV  NOT_2934(g5734,I9290);
  IV  NOT_2935(g10819,I16525);
  IV  NOT_2936(g11428,I17337);
  IV  NOT_2937(g10910,I16682);
  IV  NOT_2938(g3290,I6461);
  IV  NOT_2939(I17362,g11376);
  IV  NOT_2940(g10202,g10171);
  IV  NOT_2941(I10334,g6003);
  IV  NOT_2942(g10257,g10197);
  IV  NOT_2943(g4317,I7586);
  IV  NOT_2944(g8278,I13206);
  IV  NOT_2945(I4876,g580);
  IV  NOT_2946(g3093,I6299);
  IV  NOT_2947(g1998,g802);
  IV  NOT_2948(g5474,I8889);
  IV  NOT_2949(g10111,I15347);
  IV  NOT_2950(g7192,g6742);
  IV  NOT_2951(g5992,I9608);
  IV  NOT_2952(g7085,I11318);
  IV  NOT_2953(g3256,I6424);
  IV  NOT_2954(I7746,g3763);
  IV  NOT_2955(g6634,I10589);
  IV  NOT_2956(I9188,g4908);
  IV  NOT_2957(I10762,g6127);
  IV  NOT_2958(g8667,I13952);
  IV  NOT_2959(g3816,g3228);
  IV  NOT_2960(g8143,g8029);
  IV  NOT_2961(I13816,g8559);
  IV  NOT_2962(I15548,g10083);
  IV  NOT_2963(I6504,g3214);
  IV  NOT_2964(I9388,g5576);
  IV  NOT_2965(g8235,g7967);
  IV  NOT_2966(g8343,I13409);
  IV  NOT_2967(g6742,g5830);
  IV  NOT_2968(g11548,g11519);
  IV  NOT_2969(g6104,I9769);
  IV  NOT_2970(I14964,g9762);
  IV  NOT_2971(g10590,I16255);
  IV  NOT_2972(I9216,g4935);
  IV  NOT_2973(I6385,g2260);
  IV  NOT_2974(g6304,I10171);
  IV  NOT_2975(I16856,g10909);
  IV  NOT_2976(g8566,I13791);
  IV  NOT_2977(g6499,g5867);
  IV  NOT_2978(I16261,g10556);
  IV  NOT_2979(g2202,g148);
  IV  NOT_2980(g11504,I17531);
  IV  NOT_2981(g8988,I14385);
  IV  NOT_2982(g4775,I8139);
  IV  NOT_2983(I11752,g7032);
  IV  NOT_2984(g8134,I13005);
  IV  NOT_2985(g7941,g7406);
  IV  NOT_2986(I15317,g10025);
  IV  NOT_2987(I6025,g2259);
  IV  NOT_2988(g2908,I6077);
  IV  NOT_2989(g8334,I13382);
  IV  NOT_2990(g9265,g8892);
  IV  NOT_2991(g6926,I11046);
  IV  NOT_2992(g2094,I4924);
  IV  NOT_2993(I12415,g7631);
  IV  NOT_2994(g11317,I17112);
  IV  NOT_2995(g10094,I15329);
  IV  NOT_2996(g3397,g2896);
  IV  NOT_2997(g8548,g8390);
  IV  NOT_2998(g2518,g590);
  IV  NOT_2999(g4060,g3144);
  IV  NOT_3000(g4460,g3820);
  IV  NOT_3001(I9564,g5109);
  IV  NOT_3002(I7468,g3697);
  IV  NOT_3003(g6273,I10078);
  IV  NOT_3004(I8885,g4548);
  IV  NOT_3005(g8804,I14133);
  IV  NOT_3006(I14543,g9311);
  IV  NOT_3007(I8414,g4293);
  IV  NOT_3008(g10150,I15448);
  IV  NOT_3009(g10801,I16507);
  IV  NOT_3010(I9826,g5390);
  IV  NOT_3011(I10117,g6241);
  IV  NOT_3012(g7708,I12339);
  IV  NOT_3013(I13669,g8294);
  IV  NOT_3014(g10735,I16416);
  IV  NOT_3015(g10877,I16601);
  IV  NOT_3016(g11057,g10937);
  IV  NOT_3017(g7520,I11898);
  IV  NOT_3018(g8792,I14105);
  IV  NOT_3019(I17347,g11373);
  IV  NOT_3020(I7677,g3735);
  IV  NOT_3021(I11668,g7043);
  IV  NOT_3022(g6044,I9665);
  IV  NOT_3023(g2593,g1973);
  IV  NOT_3024(g7031,g6413);
  IV  NOT_3025(g4739,g4117);
  IV  NOT_3026(I8903,g4561);
  IV  NOT_3027(g6444,g6158);
  IV  NOT_3028(g11245,g11112);
  IV  NOT_3029(g7431,I11821);
  IV  NOT_3030(I15323,g10019);
  IV  NOT_3031(g6269,I10066);
  IV  NOT_3032(I15299,g9995);
  IV  NOT_3033(g7812,I12601);
  IV  NOT_3034(g11626,I17692);
  IV  NOT_3035(g9770,g9432);
  IV  NOT_3036(g10196,I15562);
  IV  NOT_3037(I11489,g6569);
  IV  NOT_3038(g10695,I16366);
  IV  NOT_3039(g5688,I9213);
  IV  NOT_3040(g11323,I17124);
  IV  NOT_3041(I13489,g8233);
  IV  NOT_3042(g2965,I6196);
  IV  NOT_3043(I6406,g2339);
  IV  NOT_3044(I5475,g1289);
  IV  NOT_3045(I7716,g3751);
  IV  NOT_3046(g6572,g5805);
  IV  NOT_3047(g6862,g6720);
  IV  NOT_3048(g7376,I11756);
  IV  NOT_3049(I5949,g2540);
  IV  NOT_3050(g10526,g10460);
  IV  NOT_3051(g8313,I13323);
  IV  NOT_3052(I12484,g7580);
  IV  NOT_3053(I14242,g8787);
  IV  NOT_3054(I9108,g5593);
  IV  NOT_3055(I15775,g10253);
  IV  NOT_3056(I13424,g8200);
  IV  NOT_3057(g4479,I7858);
  IV  NOT_3058(g9532,I14681);
  IV  NOT_3059(I9308,g5494);
  IV  NOT_3060(g6712,g5984);
  IV  NOT_3061(I8036,g3820);
  IV  NOT_3062(g4294,g3664);
  IV  NOT_3063(I10123,g5676);
  IV  NOT_3064(g6543,g5888);
  IV  NOT_3065(g4840,I8199);
  IV  NOT_3066(I8436,g4462);
  IV  NOT_3067(g9553,I14694);
  IV  NOT_3068(I5292,g76);
  IV  NOT_3069(I9883,g5557);
  IV  NOT_3070(I14123,g8767);
  IV  NOT_3071(g3723,g3071);
  IV  NOT_3072(g7765,I12460);
  IV  NOT_3073(g7286,I11534);
  IV  NOT_3074(g4190,I7387);
  IV  NOT_3075(I5998,g2197);
  IV  NOT_3076(g4390,g3914);
  IV  NOT_3077(I10807,g6396);
  IV  NOT_3078(g10457,I15962);
  IV  NOT_3079(g3817,I7043);
  IV  NOT_3080(g7911,g7664);
  IV  NOT_3081(I5646,g940);
  IV  NOT_3082(I10974,g6563);
  IV  NOT_3083(g8094,g7987);
  IV  NOT_3084(g2050,g1861);
  IV  NOT_3085(g2641,g1987);
  IV  NOT_3086(I8831,g4480);
  IV  NOT_3087(I15232,g9974);
  IV  NOT_3088(I10639,g5830);
  IV  NOT_3089(I17516,g11483);
  IV  NOT_3090(g2450,g1351);
  IV  NOT_3091(I16432,g10702);
  IV  NOT_3092(g4501,g3946);
  IV  NOT_3093(g8518,I13723);
  IV  NOT_3094(g6729,I10724);
  IV  NOT_3095(g6961,I11115);
  IV  NOT_3096(g8567,I13794);
  IV  NOT_3097(I10293,g5863);
  IV  NOT_3098(g4156,I7295);
  IV  NOT_3099(I11713,g7023);
  IV  NOT_3100(g7733,I12380);
  IV  NOT_3101(I5850,g2273);
  IV  NOT_3102(g7270,I11515);
  IV  NOT_3103(g9990,I15190);
  IV  NOT_3104(g6927,I11049);
  IV  NOT_3105(g3751,I6944);
  IV  NOT_3106(I9165,g5037);
  IV  NOT_3107(I16461,g10735);
  IV  NOT_3108(I9571,g5509);
  IV  NOT_3109(I9365,g5392);
  IV  NOT_3110(g7610,I12180);
  IV  NOT_3111(g2179,g89);
  IV  NOT_3112(g4942,I8308);
  IV  NOT_3113(g9029,I14424);
  IV  NOT_3114(g6014,g5309);
  IV  NOT_3115(g7073,I11296);
  IV  NOT_3116(I12799,g7556);
  IV  NOT_3117(g7796,I12553);
  IV  NOT_3118(I12813,g7688);
  IV  NOT_3119(g6885,I10979);
  IV  NOT_3120(g9429,g9082);
  IV  NOT_3121(g22,I4777);
  IV  NOT_3122(g7473,g7148);
  IV  NOT_3123(I10391,g5838);
  IV  NOT_3124(I17209,g11289);
  IV  NOT_3125(g6660,I10623);
  IV  NOT_3126(I11255,g6547);
  IV  NOT_3127(g10256,g10140);
  IV  NOT_3128(I6173,g2125);
  IV  NOT_3129(g11512,I17555);
  IV  NOT_3130(I13255,g8270);
  IV  NOT_3131(I14391,g8928);
  IV  NOT_3132(I16650,g10776);
  IV  NOT_3133(I6373,g2024);
  IV  NOT_3134(I6091,g2270);
  IV  NOT_3135(g5183,g4640);
  IV  NOT_3136(g7124,I11363);
  IV  NOT_3137(g7980,I12786);
  IV  NOT_3138(g7324,I11620);
  IV  NOT_3139(g10280,g10160);
  IV  NOT_3140(g6903,I11005);
  IV  NOT_3141(g2777,g2276);
  IV  NOT_3142(I5919,g2530);
  IV  NOT_3143(I11188,g6513);
  IV  NOT_3144(g7069,I11286);
  IV  NOT_3145(I12805,g7684);
  IV  NOT_3146(I13188,g8171);
  IV  NOT_3147(g5779,I9371);
  IV  NOT_3148(I13678,g8306);
  IV  NOT_3149(I14579,g9272);
  IV  NOT_3150(g4954,g4509);
  IV  NOT_3151(g4250,g3698);
  IV  NOT_3152(g4163,I7308);
  IV  NOT_3153(I5952,g2506);
  IV  NOT_3154(g2882,I6034);
  IV  NOT_3155(g7540,I11956);
  IV  NOT_3156(g8160,I13057);
  IV  NOT_3157(g4363,I7654);
  IV  NOT_3158(I11686,g7039);
  IV  NOT_3159(I16528,g10732);
  IV  NOT_3160(I7577,g4124);
  IV  NOT_3161(I5276,g1411);
  IV  NOT_3162(g8360,I13460);
  IV  NOT_3163(I16843,g10898);
  IV  NOT_3164(I6007,g2199);
  IV  NOT_3165(g5423,g4300);
  IV  NOT_3166(I13460,g8155);
  IV  NOT_3167(I17453,g11451);
  IV  NOT_3168(I11383,g6385);
  IV  NOT_3169(g2271,g877);
  IV  NOT_3170(g7377,I11759);
  IV  NOT_3171(g7206,I11436);
  IV  NOT_3172(g10157,I15467);
  IV  NOT_3173(g11445,I17384);
  IV  NOT_3174(g6036,I9647);
  IV  NOT_3175(I5561,g869);
  IV  NOT_3176(I13030,g8052);
  IV  NOT_3177(g2611,I5734);
  IV  NOT_3178(g4453,I7810);
  IV  NOT_3179(g8450,I13648);
  IV  NOT_3180(g6178,g4977);
  IV  NOT_3181(I6767,g2914);
  IV  NOT_3182(g11499,I17516);
  IV  NOT_3183(I8495,g4325);
  IV  NOT_3184(g3368,g3138);
  IV  NOT_3185(g9745,g9454);
  IV  NOT_3186(I11065,g6750);
  IV  NOT_3187(I6535,g2826);
  IV  NOT_3188(g1987,g762);
  IV  NOT_3189(g9338,I14519);
  IV  NOT_3190(g7287,I11537);
  IV  NOT_3191(g2799,g2276);
  IV  NOT_3192(g11498,I17513);
  IV  NOT_3193(I5986,g2194);
  IV  NOT_3194(g6135,I9842);
  IV  NOT_3195(g5665,I9156);
  IV  NOT_3196(g9109,I14452);
  IV  NOT_3197(g6335,I10228);
  IV  NOT_3198(I15989,g10417);
  IV  NOT_3199(g9309,g8892);
  IV  NOT_3200(g3531,g2971);
  IV  NOT_3201(I8869,g4421);
  IV  NOT_3202(g5127,I8535);
  IV  NOT_3203(g3458,g3144);
  IV  NOT_3204(g6182,g5446);
  IV  NOT_3205(g6288,I10123);
  IV  NOT_3206(I17274,g11389);
  IV  NOT_3207(g6382,I10278);
  IV  NOT_3208(I9662,g5319);
  IV  NOT_3209(g8179,I13086);
  IV  NOT_3210(g7849,I12644);
  IV  NOT_3211(g10876,I16598);
  IV  NOT_3212(g10885,g10809);
  IV  NOT_3213(g11056,g10950);
  IV  NOT_3214(g3743,I6932);
  IV  NOT_3215(g8379,I13485);
  IV  NOT_3216(g4912,I8282);
  IV  NOT_3217(I14116,g8766);
  IV  NOT_3218(g2997,g2135);
  IV  NOT_3219(g11611,I17657);
  IV  NOT_3220(I12400,g7537);
  IV  NOT_3221(g2541,I5658);
  IV  NOT_3222(g11080,I16853);
  IV  NOT_3223(I7426,g3334);
  IV  NOT_3224(I9290,g5052);
  IV  NOT_3225(g5146,g4596);
  IV  NOT_3226(g10854,g10708);
  IV  NOT_3227(g6805,I10825);
  IV  NOT_3228(g5633,g4388);
  IV  NOT_3229(g3505,I6694);
  IV  NOT_3230(g7781,I12508);
  IV  NOT_3231(I5970,g2185);
  IV  NOT_3232(g6749,I10756);
  IV  NOT_3233(I16708,g10822);
  IV  NOT_3234(g2238,I5237);
  IV  NOT_3235(g11432,I17347);
  IV  NOT_3236(I13837,g8488);
  IV  NOT_3237(g3411,I6616);
  IV  NOT_3238(I9093,g5397);
  IV  NOT_3239(g7900,g7712);
  IV  NOT_3240(I16258,g10555);
  IV  NOT_3241(I4948,g586);
  IV  NOT_3242(g2209,g93);
  IV  NOT_3243(g7797,I12556);
  IV  NOT_3244(I9256,g5078);
  IV  NOT_3245(I8265,g4602);
  IV  NOT_3246(I9816,g5576);
  IV  NOT_3247(g5696,I9229);
  IV  NOT_3248(I15461,g10074);
  IV  NOT_3249(g6947,I11085);
  IV  NOT_3250(I7984,g3621);
  IV  NOT_3251(I5224,g61);
  IV  NOT_3252(I7280,g3208);
  IV  NOT_3253(I10237,g6120);
  IV  NOT_3254(g6798,I10804);
  IV  NOT_3255(I8442,g4464);
  IV  NOT_3256(I12538,g7658);
  IV  NOT_3257(g8271,I13185);
  IV  NOT_3258(g2802,g2276);
  IV  NOT_3259(g11342,I17149);
  IV  NOT_3260(I10340,g6205);
  IV  NOT_3261(g1991,g778);
  IV  NOT_3262(I5120,g622);
  IV  NOT_3263(g3474,I6679);
  IV  NOT_3264(g9449,g9094);
  IV  NOT_3265(g6560,g5759);
  IV  NOT_3266(I14340,g8820);
  IV  NOT_3267(g5753,I9329);
  IV  NOT_3268(I8164,g3566);
  IV  NOT_3269(I15736,g10258);
  IV  NOT_3270(g10456,I15959);
  IV  NOT_3271(g5508,I8929);
  IV  NOT_3272(g11199,g11112);
  IV  NOT_3273(I14684,g9124);
  IV  NOT_3274(g11650,I17752);
  IV  NOT_3275(g7144,I11387);
  IV  NOT_3276(I11617,g6839);
  IV  NOT_3277(g7344,I11680);
  IV  NOT_3278(g5072,I8442);
  IV  NOT_3279(I7636,g3330);
  IV  NOT_3280(I13915,g8451);
  IV  NOT_3281(g5472,I8885);
  IV  NOT_3282(g8981,I14364);
  IV  NOT_3283(I9421,g5063);
  IV  NOT_3284(g8674,I13959);
  IV  NOT_3285(I5789,g2162);
  IV  NOT_3286(g5043,g4840);
  IV  NOT_3287(I11201,g6522);
  IV  NOT_3288(g10314,I15744);
  IV  NOT_3289(g7259,I11494);
  IV  NOT_3290(g5443,I8872);
  IV  NOT_3291(g6208,I9953);
  IV  NOT_3292(I7790,g3782);
  IV  NOT_3293(I16879,g10936);
  IV  NOT_3294(g6302,I10165);
  IV  NOT_3295(g10307,I15729);
  IV  NOT_3296(I15365,g10025);
  IV  NOT_3297(I7061,g3050);
  IV  NOT_3298(g6579,g5949);
  IV  NOT_3299(g5116,g4682);
  IV  NOT_3300(g6869,I10949);
  IV  NOT_3301(g7852,g7479);
  IV  NOT_3302(g7923,g7527);
  IV  NOT_3303(I17164,g11320);
  IV  NOT_3304(I7387,g4083);
  IV  NOT_3305(g10596,I16269);
  IV  NOT_3306(I11467,g6488);
  IV  NOT_3307(I11494,g6574);
  IV  NOT_3308(I13595,g8339);
  IV  NOT_3309(g8132,I12999);
  IV  NOT_3310(g6719,I10710);
  IV  NOT_3311(I12235,g7082);
  IV  NOT_3312(g8332,I13376);
  IV  NOT_3313(g10243,I15635);
  IV  NOT_3314(I11623,g6841);
  IV  NOT_3315(I12683,g7387);
  IV  NOT_3316(I6388,g2329);
  IV  NOT_3317(g8680,I13965);
  IV  NOT_3318(g10431,g10328);
  IV  NOT_3319(I11037,g6629);
  IV  NOT_3320(g8353,I13439);
  IV  NOT_3321(I14130,g8769);
  IV  NOT_3322(I10362,g6224);
  IV  NOT_3323(g2864,g2298);
  IV  NOT_3324(I10165,g5948);
  IV  NOT_3325(I13782,g8515);
  IV  NOT_3326(g6917,I11029);
  IV  NOT_3327(g4894,I8247);
  IV  NOT_3328(I6028,g2208);
  IV  NOT_3329(g10269,g10154);
  IV  NOT_3330(g8802,I14127);
  IV  NOT_3331(I6671,g2757);
  IV  NOT_3332(I6428,g2348);
  IV  NOT_3333(g7886,g7479);
  IV  NOT_3334(g4735,g3546);
  IV  NOT_3335(I17327,g11349);
  IV  NOT_3336(g6265,I10054);
  IV  NOT_3337(g3976,I7109);
  IV  NOT_3338(I6247,g2462);
  IV  NOT_3339(g4782,g4089);
  IV  NOT_3340(I11155,g6470);
  IV  NOT_3341(g10156,I15464);
  IV  NOT_3342(I15708,g10241);
  IV  NOT_3343(I17537,g11497);
  IV  NOT_3344(I13418,g8145);
  IV  NOT_3345(I13822,g8488);
  IV  NOT_3346(g5697,I9232);
  IV  NOT_3347(I10006,g5633);
  IV  NOT_3348(g6442,I10362);
  IV  NOT_3349(g9452,I14645);
  IV  NOT_3350(g7314,I11590);
  IV  NOT_3351(g5210,I8631);
  IV  NOT_3352(I17108,g11225);
  IV  NOT_3353(g11471,I17450);
  IV  NOT_3354(I7345,g4050);
  IV  NOT_3355(I16458,g10734);
  IV  NOT_3356(I8429,g4458);
  IV  NOT_3357(I9605,g5620);
  IV  NOT_3358(g4475,I7852);
  IV  NOT_3359(g5596,I9020);
  IV  NOT_3360(g6164,g5426);
  IV  NOT_3361(I7763,g3769);
  IV  NOT_3362(I7191,g2646);
  IV  NOT_3363(g10734,I16413);
  IV  NOT_3364(I10437,g5755);
  IV  NOT_3365(g10335,I15787);
  IV  NOT_3366(g7650,I12261);
  IV  NOT_3367(g3326,I6495);
  IV  NOT_3368(I15244,g10031);
  IV  NOT_3369(g4292,g3863);
  IV  NOT_3370(g10930,g10827);
  IV  NOT_3371(g11043,I16790);
  IV  NOT_3372(g6454,I10388);
  IV  NOT_3373(g11244,g11112);
  IV  NOT_3374(g4526,I7931);
  IV  NOT_3375(I5478,g1212);
  IV  NOT_3376(g6296,I10147);
  IV  NOT_3377(I11194,g6515);
  IV  NOT_3378(g3760,g3003);
  IV  NOT_3379(g7008,I11149);
  IV  NOT_3380(I13194,g8140);
  IV  NOT_3381(I13589,g8361);
  IV  NOT_3382(g2623,g1999);
  IV  NOT_3383(I17381,g11436);
  IV  NOT_3384(I7536,g4098);
  IV  NOT_3385(I9585,g5241);
  IV  NOT_3386(g2076,I4886);
  IV  NOT_3387(g10131,I15395);
  IV  NOT_3388(g2889,I6049);
  IV  NOT_3389(I11524,g6593);
  IV  NOT_3390(I16598,g10804);
  IV  NOT_3391(g11069,g10974);
  IV  NOT_3392(g4084,g3119);
  IV  NOT_3393(I11836,g7220);
  IV  NOT_3394(I5435,g18);
  IV  NOT_3395(g4603,g3829);
  IV  NOT_3396(g5936,I9564);
  IV  NOT_3397(g7336,I11656);
  IV  NOT_3398(g8600,g8475);
  IV  NOT_3399(I15068,g9710);
  IV  NOT_3400(g7768,I12469);
  IV  NOT_3401(g4439,I7793);
  IV  NOT_3402(g11657,I17773);
  IV  NOT_3403(g5117,g4682);
  IV  NOT_3404(g6553,I10477);
  IV  NOT_3405(g8714,I14005);
  IV  NOT_3406(g11068,g10974);
  IV  NOT_3407(I7858,g3631);
  IV  NOT_3408(I11477,g6488);
  IV  NOT_3409(g7594,I12120);
  IV  NOT_3410(g10487,I16098);
  IV  NOT_3411(g7972,I12770);
  IV  NOT_3412(g2175,g44);
  IV  NOT_3413(I11119,g6461);
  IV  NOT_3414(g9025,I14412);
  IV  NOT_3415(g2871,I6013);
  IV  NOT_3416(g10619,I16292);
  IV  NOT_3417(I12759,g7702);
  IV  NOT_3418(I7757,g3767);
  IV  NOT_3419(I16817,g10912);
  IV  NOT_3420(I9673,g5182);
  IV  NOT_3421(I14236,g8802);
  IV  NOT_3422(g7806,I12583);
  IV  NOT_3423(I10952,g6556);
  IV  NOT_3424(g3220,I6398);
  IV  NOT_3425(I8109,g3622);
  IV  NOT_3426(g2651,g2007);
  IV  NOT_3427(I6217,g2302);
  IV  NOT_3428(g4583,g3880);
  IV  NOT_3429(g6412,I10322);
  IV  NOT_3430(I17390,g11430);
  IV  NOT_3431(g10279,g10158);
  IV  NOT_3432(g7065,I11272);
  IV  NOT_3433(I7315,g2891);
  IV  NOT_3434(g6389,I10289);
  IV  NOT_3435(I7642,g3440);
  IV  NOT_3436(I9168,g5040);
  IV  NOT_3437(g6706,I10685);
  IV  NOT_3438(I9669,g5426);
  IV  NOT_3439(g7887,g7693);
  IV  NOT_3440(g7122,I11357);
  IV  NOT_3441(I15792,g10279);
  IV  NOT_3442(I9368,g5288);
  IV  NOT_3443(g7322,I11614);
  IV  NOT_3444(g4919,I8290);
  IV  NOT_3445(I10063,g5766);
  IV  NOT_3446(g6990,I11132);
  IV  NOT_3447(I7447,g3694);
  IV  NOT_3448(g10278,g10182);
  IV  NOT_3449(g3977,I7112);
  IV  NOT_3450(I6861,g2942);
  IV  NOT_3451(g6888,I10984);
  IV  NOT_3452(I16656,g10791);
  IV  NOT_3453(I9531,g5004);
  IV  NOT_3454(g6171,g5446);
  IV  NOT_3455(g2184,g1806);
  IV  NOT_3456(I16295,g10552);
  IV  NOT_3457(I9458,g5091);
  IV  NOT_3458(g3161,I6367);
  IV  NOT_3459(I11704,g7008);
  IV  NOT_3460(I12849,g7632);
  IV  NOT_3461(I6055,g2569);
  IV  NOT_3462(I17522,g11485);
  IV  NOT_3463(g2339,I5399);
  IV  NOT_3464(g7033,I11188);
  IV  NOT_3465(g10039,I15244);
  IV  NOT_3466(I10873,g6331);
  IV  NOT_3467(g6956,I11106);
  IV  NOT_3468(g5597,I9023);
  IV  NOT_3469(I14873,g9525);
  IV  NOT_3470(I7654,g3728);
  IV  NOT_3471(I13809,g8480);
  IV  NOT_3472(I6133,g2253);
  IV  NOT_3473(g3051,g2135);
  IV  NOT_3474(g2838,g2165);
  IV  NOT_3475(g8076,I12930);
  IV  NOT_3476(g2024,g1718);
  IV  NOT_3477(I15458,g10069);
  IV  NOT_3478(I13466,g8160);
  IV  NOT_3479(I9505,g5088);
  IV  NOT_3480(g6281,I10102);
  IV  NOT_3481(g8476,I13674);
  IV  NOT_3482(g3327,I6498);
  IV  NOT_3483(g2424,g1690);
  IV  NOT_3484(I8449,g4469);
  IV  NOT_3485(I12652,g7458);
  IV  NOT_3486(g9766,g9432);
  IV  NOT_3487(g2809,I5909);
  IV  NOT_3488(g5784,I9380);
  IV  NOT_3489(g4004,I7140);
  IV  NOT_3490(I9734,g5257);
  IV  NOT_3491(I13036,g8053);
  IV  NOT_3492(I5002,g1173);
  IV  NOT_3493(I8865,g4518);
  IV  NOT_3494(g7550,g6974);
  IV  NOT_3495(g6297,I10150);
  IV  NOT_3496(I11560,g7037);
  IV  NOT_3497(g10187,I15539);
  IV  NOT_3498(I6196,g2462);
  IV  NOT_3499(I5824,g2502);
  IV  NOT_3500(g7845,I12634);
  IV  NOT_3501(I10834,g6715);
  IV  NOT_3502(g8871,I14185);
  IV  NOT_3503(g8375,I13475);
  IV  NOT_3504(I15545,g10075);
  IV  NOT_3505(g3633,I6802);
  IV  NOT_3506(I15079,g9745);
  IV  NOT_3507(I8098,g3583);
  IV  NOT_3508(g2077,g219);
  IV  NOT_3509(g2231,I5218);
  IV  NOT_3510(g7195,I11417);
  IV  NOT_3511(g11545,g11519);
  IV  NOT_3512(g11079,I16850);
  IV  NOT_3513(g11444,I17381);
  IV  NOT_3514(g5937,I9567);
  IV  NOT_3515(g7395,g6941);
  IV  NOT_3516(I13642,g8378);
  IV  NOT_3517(g7337,I11659);
  IV  NOT_3518(g3103,g2391);
  IV  NOT_3519(I9074,g4764);
  IV  NOT_3520(g7913,g7467);
  IV  NOT_3521(I6538,g2827);
  IV  NOT_3522(g2523,I5632);
  IV  NOT_3523(I7272,g3253);
  IV  NOT_3524(g2643,g1989);
  IV  NOT_3525(I9992,g5633);
  IV  NOT_3526(g10143,I15427);
  IV  NOT_3527(g5668,I9165);
  IV  NOT_3528(g11078,I16847);
  IV  NOT_3529(g6338,I10237);
  IV  NOT_3530(I15598,g10170);
  IV  NOT_3531(I10021,g5692);
  IV  NOT_3532(g5840,g5320);
  IV  NOT_3533(g4970,g4411);
  IV  NOT_3534(g8500,I13695);
  IV  NOT_3535(I7612,g3817);
  IV  NOT_3536(g11598,I17642);
  IV  NOT_3537(I7017,g3068);
  IV  NOT_3538(g6109,g5052);
  IV  NOT_3539(I12406,g7464);
  IV  NOT_3540(g6309,I10186);
  IV  NOT_3541(g11086,I16867);
  IV  NOT_3542(g7807,I12586);
  IV  NOT_3543(I7417,g4160);
  IV  NOT_3544(g3732,I6914);
  IV  NOT_3545(I17252,g11343);
  IV  NOT_3546(g10169,I15503);
  IV  NOT_3547(I7935,g3440);
  IV  NOT_3548(I9080,g4775);
  IV  NOT_3549(g8184,I13105);
  IV  NOT_3550(g10884,g10809);
  IV  NOT_3551(g6808,I10834);
  IV  NOT_3552(I15817,g10199);
  IV  NOT_3553(I9863,g5557);
  IV  NOT_3554(g8139,g8025);
  IV  NOT_3555(I16289,g10541);
  IV  NOT_3556(g8339,I13397);
  IV  NOT_3557(g2742,I5798);
  IV  NOT_3558(g3944,g2920);
  IV  NOT_3559(g10168,I15500);
  IV  NOT_3560(I10607,g5763);
  IV  NOT_3561(g6707,g5949);
  IV  NOT_3562(I13630,g8334);
  IV  NOT_3563(g2304,I5348);
  IV  NOT_3564(g11322,I17121);
  IV  NOT_3565(g9091,g8892);
  IV  NOT_3566(g4320,g4013);
  IV  NOT_3567(I15977,g10411);
  IV  NOT_3568(g11159,g10950);
  IV  NOT_3569(I10274,g5811);
  IV  NOT_3570(I11166,g6480);
  IV  NOT_3571(I11665,g7038);
  IV  NOT_3572(I16571,g10819);
  IV  NOT_3573(I13166,g8009);
  IV  NOT_3574(I7330,g3761);
  IV  NOT_3575(I8268,g4674);
  IV  NOT_3576(g8424,I13586);
  IV  NOT_3577(I5064,g1690);
  IV  NOT_3578(g8795,I14112);
  IV  NOT_3579(g10217,I15589);
  IV  NOT_3580(g7142,I11383);
  IV  NOT_3581(I6256,g2462);
  IV  NOT_3582(g4277,g3688);
  IV  NOT_3583(g6201,I9938);
  IV  NOT_3584(g7342,I11674);
  IV  NOT_3585(I11008,g6795);
  IV  NOT_3586(g6957,I11109);
  IV  NOT_3587(I15353,g10007);
  IV  NOT_3588(g2754,I5830);
  IV  NOT_3589(g4906,I8275);
  IV  NOT_3590(g7815,I12610);
  IV  NOT_3591(g11656,I17770);
  IV  NOT_3592(g4789,g3337);
  IV  NOT_3593(I7800,g3791);
  IV  NOT_3594(g10486,I16095);
  IV  NOT_3595(g11353,I17176);
  IV  NOT_3596(g8077,I12933);
  IV  NOT_3597(I15823,g10201);
  IV  NOT_3598(g6449,g6172);
  IV  NOT_3599(I13485,g8194);
  IV  NOT_3600(g2273,g881);
  IV  NOT_3601(g8477,g8317);
  IV  NOT_3602(g6575,g5949);
  IV  NOT_3603(g7692,g7148);
  IV  NOT_3604(I12613,g7525);
  IV  NOT_3605(g8523,I13732);
  IV  NOT_3606(I6381,g2257);
  IV  NOT_3607(g9767,I14914);
  IV  NOT_3608(g7097,I11330);
  IV  NOT_3609(I9688,g5201);
  IV  NOT_3610(g7726,I12363);
  IV  NOT_3611(I9857,g5269);
  IV  NOT_3612(I13454,g8183);
  IV  NOT_3613(g2613,I5740);
  IV  NOT_3614(g7497,g7148);
  IV  NOT_3615(g9535,I14690);
  IV  NOT_3616(g6715,I10702);
  IV  NOT_3617(g2044,I4850);
  IV  NOT_3618(g7354,I11710);
  IV  NOT_3619(g10580,g10530);
  IV  NOT_3620(I10153,g5947);
  IV  NOT_3621(g2444,g876);
  IV  NOT_3622(I5237,g1107);
  IV  NOT_3623(g5032,I8403);
  IV  NOT_3624(g2269,I5308);
  IV  NOT_3625(g10223,I15595);
  IV  NOT_3626(I7213,g2635);
  IV  NOT_3627(g9261,g8892);
  IV  NOT_3628(I6421,g2346);
  IV  NOT_3629(g4299,g4144);
  IV  NOT_3630(I14409,g8938);
  IV  NOT_3631(I12463,g7579);
  IV  NOT_3632(g3697,I6856);
  IV  NOT_3633(g8099,g7990);
  IV  NOT_3634(I8385,g4238);
  IV  NOT_3635(I14136,g8775);
  IV  NOT_3636(g8304,I13280);
  IV  NOT_3637(g3914,g3015);
  IV  NOT_3638(I9126,g4891);
  IV  NOT_3639(I13239,g8266);
  IV  NOT_3640(g10110,I15344);
  IV  NOT_3641(g11631,I17707);
  IV  NOT_3642(I9326,g5320);
  IV  NOT_3643(g2543,I5662);
  IV  NOT_3644(g6584,I10538);
  IV  NOT_3645(g11017,I16742);
  IV  NOT_3646(g6539,I10461);
  IV  NOT_3647(g6896,I10996);
  IV  NOT_3648(g5568,I8985);
  IV  NOT_3649(g10321,I15759);
  IV  NOT_3650(I5089,g1854);
  IV  NOT_3651(I5731,g2089);
  IV  NOT_3652(I11238,g6543);
  IV  NOT_3653(I17213,g11290);
  IV  NOT_3654(g7783,I12514);
  IV  NOT_3655(g10179,g10041);
  IV  NOT_3656(g10531,g10471);
  IV  NOT_3657(g7979,I12783);
  IV  NOT_3658(g3413,g2896);
  IV  NOT_3659(g5912,I9544);
  IV  NOT_3660(g7312,I11584);
  IV  NOT_3661(I7166,g2620);
  IV  NOT_3662(I5966,g2541);
  IV  NOT_3663(g10178,I15526);
  IV  NOT_3664(I7366,g4012);
  IV  NOT_3665(g4738,g3440);
  IV  NOT_3666(I13941,g8488);
  IV  NOT_3667(I13382,g8134);
  IV  NOT_3668(g6268,I10063);
  IV  NOT_3669(I11519,g6591);
  IV  NOT_3670(I11176,g6501);
  IV  NOT_3671(g10186,I15536);
  IV  NOT_3672(g7001,I11140);
  IV  NOT_3673(g8273,I13191);
  IV  NOT_3674(g10676,g10570);
  IV  NOT_3675(g6419,I10331);
  IV  NOT_3676(I10891,g6334);
  IV  NOT_3677(I13185,g8192);
  IV  NOT_3678(g11289,I17070);
  IV  NOT_3679(I7456,g3716);
  IV  NOT_3680(g1993,g786);
  IV  NOT_3681(g3820,I7048);
  IV  NOT_3682(g7676,I12303);
  IV  NOT_3683(g4140,I7284);
  IV  NOT_3684(g6052,g5426);
  IV  NOT_3685(g11309,I17096);
  IV  NOT_3686(g4078,I7205);
  IV  NOT_3687(I12514,g7735);
  IV  NOT_3688(g8613,g8484);
  IV  NOT_3689(I16525,g10719);
  IV  NOT_3690(I7348,g4056);
  IV  NOT_3691(g6452,I10384);
  IV  NOT_3692(I9383,g5296);
  IV  NOT_3693(I9608,g5127);
  IV  NOT_3694(I15308,g10019);
  IV  NOT_3695(g7329,I11635);
  IV  NOT_3696(g4478,g3820);
  IV  NOT_3697(g7761,I12448);
  IV  NOT_3698(g2014,g1104);
  IV  NOT_3699(g4907,I8278);
  IV  NOT_3700(g8444,I13630);
  IV  NOT_3701(g2885,I6043);
  IV  NOT_3702(I9779,g5391);
  IV  NOT_3703(g2946,I6133);
  IV  NOT_3704(g4435,g3914);
  IV  NOT_3705(I9023,g4727);
  IV  NOT_3706(g8983,I14370);
  IV  NOT_3707(g4082,I7213);
  IV  NOT_3708(I12421,g7634);
  IV  NOT_3709(I8406,g4274);
  IV  NOT_3710(I5254,g1700);
  IV  NOT_3711(I14109,g8765);
  IV  NOT_3712(g8572,I13809);
  IV  NOT_3713(g7727,I12366);
  IV  NOT_3714(I7964,g3433);
  IV  NOT_3715(g2903,g2166);
  IV  NOT_3716(I7260,g2844);
  IV  NOT_3717(I14537,g9308);
  IV  NOT_3718(I10108,g5743);
  IV  NOT_3719(g6086,I9737);
  IV  NOT_3720(g8712,g8680);
  IV  NOT_3721(g11495,I17500);
  IV  NOT_3722(I12012,g6916);
  IV  NOT_3723(I9588,g5114);
  IV  NOT_3724(g7746,I12403);
  IV  NOT_3725(I8487,g4526);
  IV  NOT_3726(I5438,g18);
  IV  NOT_3727(g3775,I7002);
  IV  NOT_3728(g7221,I11459);
  IV  NOT_3729(I17350,g11377);
  IV  NOT_3730(I14303,g8811);
  IV  NOT_3731(g6385,g6119);
  IV  NOT_3732(g6881,I10971);
  IV  NOT_3733(I12541,g7662);
  IV  NOT_3734(g7703,g7085);
  IV  NOT_3735(I9665,g5174);
  IV  NOT_3736(I15752,g10264);
  IV  NOT_3737(g4915,g4413);
  IV  NOT_3738(g2178,g45);
  IV  NOT_3739(g2436,I5525);
  IV  NOT_3740(I15374,g10007);
  IV  NOT_3741(g9028,I14421);
  IV  NOT_3742(g8729,g8595);
  IV  NOT_3743(g8961,I14330);
  IV  NOT_3744(I4900,g583);
  IV  NOT_3745(I11501,g6581);
  IV  NOT_3746(I16610,g10792);
  IV  NOT_3747(g9671,I14802);
  IV  NOT_3748(I17152,g11308);
  IV  NOT_3749(g3060,g2135);
  IV  NOT_3750(I13729,g8290);
  IV  NOT_3751(I13577,g8330);
  IV  NOT_3752(I10381,g5847);
  IV  NOT_3753(g4214,I7459);
  IV  NOT_3754(I16255,g10554);
  IV  NOT_3755(I14982,g9672);
  IV  NOT_3756(g6425,g6141);
  IV  NOT_3757(I11728,g7010);
  IV  NOT_3758(g11643,I17733);
  IV  NOT_3759(g2135,I5064);
  IV  NOT_3760(I16679,g10784);
  IV  NOT_3761(g2335,I5391);
  IV  NOT_3762(g5683,I9202);
  IV  NOT_3763(I13439,g8187);
  IV  NOT_3764(I9346,g5281);
  IV  NOT_3765(I7118,g2979);
  IV  NOT_3766(g4310,I7577);
  IV  NOT_3767(g2382,g599);
  IV  NOT_3768(I7318,g3266);
  IV  NOT_3769(I12829,g7680);
  IV  NOT_3770(I16124,g10396);
  IV  NOT_3771(g10909,I16679);
  IV  NOT_3772(I12535,g7656);
  IV  NOT_3773(g5778,I9368);
  IV  NOT_3774(I10174,g5994);
  IV  NOT_3775(I15669,g10194);
  IV  NOT_3776(g10543,I16196);
  IV  NOT_3777(g3784,g2586);
  IV  NOT_3778(I17413,g11425);
  IV  NOT_3779(g5894,g5361);
  IV  NOT_3780(g9826,I14979);
  IV  NOT_3781(g10117,I15359);
  IV  NOT_3782(g8660,I13945);
  IV  NOT_3783(g8946,I14295);
  IV  NOT_3784(g10908,I16676);
  IV  NOT_3785(g2916,I6097);
  IV  NOT_3786(I7843,g3440);
  IV  NOT_3787(g2022,g1346);
  IV  NOT_3788(g5735,I9293);
  IV  NOT_3789(I15392,g10104);
  IV  NOT_3790(g7677,g7148);
  IV  NOT_3791(g2749,I5815);
  IV  NOT_3792(g3995,g3121);
  IV  NOT_3793(g3937,I7086);
  IV  NOT_3794(I10840,g6719);
  IV  NOT_3795(g9741,I14888);
  IV  NOT_3796(g4002,g3121);
  IV  NOT_3797(I7393,g4096);
  IV  NOT_3798(I16938,g11086);
  IV  NOT_3799(I6531,g3186);
  IV  NOT_3800(I11348,g6695);
  IV  NOT_3801(I12344,g7062);
  IV  NOT_3802(I13083,g7921);
  IV  NOT_3803(g3479,g2655);
  IV  NOT_3804(g11195,g11112);
  IV  NOT_3805(g11489,I17482);
  IV  NOT_3806(g6131,g5548);
  IV  NOT_3807(g5661,I9144);
  IV  NOT_3808(g10747,I16432);
  IV  NOT_3809(I15559,g10094);
  IV  NOT_3810(g5075,g4439);
  IV  NOT_3811(g8513,I13708);
  IV  NOT_3812(I15488,g10116);
  IV  NOT_3813(I15424,g10080);
  IV  NOT_3814(g6406,I10314);
  IV  NOT_3815(g10242,I15632);
  IV  NOT_3816(I8007,g3829);
  IV  NOT_3817(g5475,I8892);
  IV  NOT_3818(g4762,I8116);
  IV  NOT_3819(g2798,g2449);
  IV  NOT_3820(g5949,I9591);
  IV  NOT_3821(g7349,I11695);
  IV  NOT_3822(I10192,g6115);
  IV  NOT_3823(g11424,I17327);
  IV  NOT_3824(I9240,g5069);
  IV  NOT_3825(g6635,I10592);
  IV  NOT_3826(I11566,g6820);
  IV  NOT_3827(g11016,I16739);
  IV  NOT_3828(g9108,I14449);
  IV  NOT_3829(g3390,g3161);
  IV  NOT_3830(g9308,I14499);
  IV  NOT_3831(g8036,I12878);
  IV  NOT_3832(g2560,I5684);
  IV  NOT_3833(g5627,g4840);
  IV  NOT_3834(g8436,I13606);
  IV  NOT_3835(g8178,I13083);
  IV  NOT_3836(g6801,I10813);
  IV  NOT_3837(g6305,I10174);
  IV  NOT_3838(I6856,g3318);
  IV  NOT_3839(g4590,I7999);
  IV  NOT_3840(g7848,I12641);
  IV  NOT_3841(g5292,g4445);
  IV  NOT_3842(I10663,g6040);
  IV  NOT_3843(g8378,I13482);
  IV  NOT_3844(g9883,I15060);
  IV  NOT_3845(I9043,g4786);
  IV  NOT_3846(g3501,g3077);
  IV  NOT_3847(I14522,g9108);
  IV  NOT_3848(I8535,g4340);
  IV  NOT_3849(I9443,g5557);
  IV  NOT_3850(g7747,I12406);
  IV  NOT_3851(g5998,I9620);
  IV  NOT_3852(g5646,I9099);
  IV  NOT_3853(g10974,I16723);
  IV  NOT_3854(g8335,I13385);
  IV  NOT_3855(g2873,I6019);
  IV  NOT_3856(g6748,I10753);
  IV  NOT_3857(g2632,g2002);
  IV  NOT_3858(I6074,g2228);
  IV  NOT_3859(g2095,g143);
  IV  NOT_3860(I11653,g6954);
  IV  NOT_3861(g2037,g1771);
  IV  NOT_3862(g8182,I13099);
  IV  NOT_3863(I4886,g257);
  IV  NOT_3864(g4222,g3638);
  IV  NOT_3865(g5603,I9029);
  IV  NOT_3866(I6474,g2297);
  IV  NOT_3867(I7625,g4164);
  IV  NOT_3868(g5039,I8418);
  IV  NOT_3869(I4951,g262);
  IV  NOT_3870(g10293,I15701);
  IV  NOT_3871(g2653,g2011);
  IV  NOT_3872(g2208,g84);
  IV  NOT_3873(g2302,g29);
  IV  NOT_3874(I12029,g6922);
  IV  NOT_3875(g5850,g5320);
  IV  NOT_3876(g6226,I9973);
  IV  NOT_3877(I10553,g6192);
  IV  NOT_3878(g3704,I6861);
  IV  NOT_3879(g8805,I14136);
  IV  NOT_3880(g10265,g10143);
  IV  NOT_3881(g2579,g1969);
  IV  NOT_3882(I5837,g2507);
  IV  NOT_3883(I7938,g3406);
  IV  NOT_3884(I9147,g5011);
  IV  NOT_3885(I13636,g8357);
  IV  NOT_3886(g8422,I13580);
  IV  NOT_3887(I10949,g6747);
  IV  NOT_3888(I17302,g11391);
  IV  NOT_3889(g4899,I8262);
  IV  NOT_3890(I11333,g6670);
  IV  NOT_3891(I13415,g8144);
  IV  NOT_3892(g4464,I7829);
  IV  NOT_3893(g2719,g2043);
  IV  NOT_3894(g9448,g9091);
  IV  NOT_3895(I7909,g3387);
  IV  NOT_3896(I6080,g2108);
  IV  NOT_3897(I14326,g8818);
  IV  NOT_3898(g4785,g3337);
  IV  NOT_3899(g11042,I16787);
  IV  NOT_3900(g10391,g10313);
  IV  NOT_3901(I6480,g2462);
  IV  NOT_3902(g5702,I9243);
  IV  NOT_3903(g6445,I10367);
  IV  NOT_3904(g2752,I5824);
  IV  NOT_3905(I14040,g8649);
  IV  NOT_3906(I14948,g9555);
  IV  NOT_3907(g9827,I14982);
  IV  NOT_3908(g6091,I9744);
  IV  NOT_3909(I10702,g6071);
  IV  NOT_3910(g3810,g3228);
  IV  NOT_3911(g3363,I6549);
  IV  NOT_3912(I10904,g6558);
  IV  NOT_3913(g8798,I14119);
  IV  NOT_3914(g7119,I11354);
  IV  NOT_3915(g7319,I11605);
  IV  NOT_3916(g3432,g3144);
  IV  NOT_3917(I6569,g3186);
  IV  NOT_3918(g10579,g10528);
  IV  NOT_3919(g4563,g3946);
  IV  NOT_3920(g9774,g9474);
  IV  NOT_3921(I7606,g4166);
  IV  NOT_3922(g8560,I13773);
  IV  NOT_3923(I14252,g8783);
  IV  NOT_3924(g6169,I9896);
  IV  NOT_3925(I15383,g10107);
  IV  NOT_3926(I16277,g10536);
  IV  NOT_3927(g6283,I10108);
  IV  NOT_3928(g7352,I11704);
  IV  NOT_3929(g2042,g1796);
  IV  NOT_3930(g4295,I7556);
  IV  NOT_3931(g10578,g10527);
  IV  NOT_3932(I9013,g4767);
  IV  NOT_3933(g4237,g4013);
  IV  NOT_3934(g6407,I10317);
  IV  NOT_3935(I14564,g9026);
  IV  NOT_3936(g6920,I11034);
  IV  NOT_3937(g6578,I10526);
  IV  NOT_3938(g6868,I10946);
  IV  NOT_3939(g5616,I9046);
  IV  NOT_3940(I16595,g10783);
  IV  NOT_3941(g8873,I14191);
  IV  NOT_3942(g8632,I13915);
  IV  NOT_3943(g8095,g7942);
  IV  NOT_3944(g2164,I5095);
  IV  NOT_3945(g6718,g5949);
  IV  NOT_3946(g2364,g611);
  IV  NOT_3947(g2233,I5224);
  IV  NOT_3948(g9780,g9474);
  IV  NOT_3949(g4194,I7399);
  IV  NOT_3950(I16623,g10858);
  IV  NOT_3951(g8437,I13609);
  IV  NOT_3952(I10183,g6108);
  IV  NOT_3953(I7586,g4127);
  IV  NOT_3954(g11065,g10974);
  IV  NOT_3955(g4394,I7729);
  IV  NOT_3956(I5192,g55);
  IV  NOT_3957(I6976,g2884);
  IV  NOT_3958(g2054,g1864);
  IV  NOT_3959(g6582,g5949);
  IV  NOT_3960(I13609,g8312);
  IV  NOT_3961(I14397,g8888);
  IV  NOT_3962(g7386,I11767);
  IV  NOT_3963(g4731,I8085);
  IV  NOT_3964(I11312,g6488);
  IV  NOT_3965(g5647,I9102);
  IV  NOT_3966(g2454,I5549);
  IV  NOT_3967(g8579,I13822);
  IV  NOT_3968(g8869,I14179);
  IV  NOT_3969(g7975,I12773);
  IV  NOT_3970(I13200,g8251);
  IV  NOT_3971(g6261,I10042);
  IV  NOT_3972(I11608,g6903);
  IV  NOT_3973(g2296,I5332);
  IV  NOT_3974(I11115,g6462);
  IV  NOT_3975(I12604,g7630);
  IV  NOT_3976(g10116,I15356);
  IV  NOT_3977(I9117,g5615);
  IV  NOT_3978(g6793,I10795);
  IV  NOT_3979(g8719,g8579);
  IV  NOT_3980(g4557,g3946);
  IV  NOT_3981(I9317,g5576);
  IV  NOT_3982(g2725,g2018);
  IV  NOT_3983(g1974,g627);
  IV  NOT_3984(I14509,g8926);
  IV  NOT_3985(g5546,I8973);
  IV  NOT_3986(g7026,I11173);
  IV  NOT_3987(I5854,g2523);
  IV  NOT_3988(I8388,g4239);
  IV  NOT_3989(g4966,I8340);
  IV  NOT_3990(I12770,g7638);
  IV  NOT_3991(I14933,g9454);
  IV  NOT_3992(g7426,I11814);
  IV  NOT_3993(g9994,I15196);
  IV  NOT_3994(g9290,I14494);
  IV  NOT_3995(I11921,g6904);
  IV  NOT_3996(I17662,g11602);
  IV  NOT_3997(I12981,g8041);
  IV  NOT_3998(g8752,g8635);
  IV  NOT_3999(g6227,g5446);
  IV  NOT_4000(g10041,I15250);
  IV  NOT_4001(g5503,g4515);
  IV  NOT_4002(I7710,g3749);
  IV  NOT_4003(g7614,I12190);
  IV  NOT_4004(g10275,I15669);
  IV  NOT_4005(g4242,g3664);
  IV  NOT_4006(g10493,I16114);
  IV  NOT_4007(g7325,I11623);
  IV  NOT_4008(I17249,g11342);
  IV  NOT_4009(g4948,I8315);
  IV  NOT_4010(I7691,g3363);
  IV  NOT_4011(g9816,g9490);
  IV  NOT_4012(I17482,g11479);
  IV  NOT_4013(g10465,I15986);
  IV  NOT_4014(g1980,g646);
  IV  NOT_4015(I8247,g4615);
  IV  NOT_4016(g7984,I12796);
  IV  NOT_4017(g2012,g981);
  IV  NOT_4018(g11160,g10950);
  IV  NOT_4019(g8442,I13624);
  IV  NOT_4020(I17710,g11620);
  IV  NOT_4021(g6203,g5446);
  IV  NOT_4022(I17552,g11502);
  IV  NOT_4023(I16853,g10907);
  IV  NOT_4024(I9581,g5111);
  IV  NOT_4025(g10035,I15241);
  IV  NOT_4026(g5120,I8520);
  IV  NOT_4027(I5031,g928);
  IV  NOT_4028(g5320,g4418);
  IV  NOT_4029(g4254,g4013);
  IV  NOT_4030(I16589,g10820);
  IV  NOT_4031(I11674,g7051);
  IV  NOT_4032(g10806,I16518);
  IV  NOT_4033(g7544,I11964);
  IV  NOT_4034(g8164,g7872);
  IV  NOT_4035(I13674,g8304);
  IV  NOT_4036(I15470,g10111);
  IV  NOT_4037(I5812,g2090);
  IV  NOT_4038(g8233,g7872);
  IV  NOT_4039(g11617,I17669);
  IV  NOT_4040(I6183,g2131);
  IV  NOT_4041(g11470,I17447);
  IV  NOT_4042(I7659,g3731);
  IV  NOT_4043(g10142,I15424);
  IV  NOT_4044(g2888,I6046);
  IV  NOT_4045(I6924,g2843);
  IV  NOT_4046(g7636,I12248);
  IV  NOT_4047(I6220,g883);
  IV  NOT_4048(I4891,g582);
  IV  NOT_4049(g2171,I5116);
  IV  NOT_4050(g4438,I7790);
  IV  NOT_4051(I14452,g8922);
  IV  NOT_4052(g4773,I8133);
  IV  NOT_4053(g7306,I11566);
  IV  NOT_4054(I13732,g8291);
  IV  NOT_4055(g8296,I13242);
  IV  NOT_4056(g2956,I6159);
  IV  NOT_4057(I15075,g9761);
  IV  NOT_4058(g8725,g8589);
  IV  NOT_4059(g7790,I12535);
  IV  NOT_4060(g9263,g8892);
  IV  NOT_4061(g3683,I6844);
  IV  NOT_4062(g11075,g10937);
  IV  NOT_4063(I5765,g2004);
  IV  NOT_4064(I15595,g10165);
  IV  NOT_4065(I15467,g10079);
  IV  NOT_4066(I15494,g10117);
  IV  NOT_4067(I17356,g11384);
  IV  NOT_4068(g8532,I13741);
  IV  NOT_4069(I8308,g4443);
  IV  NOT_4070(g7187,I11405);
  IV  NOT_4071(I7311,g2803);
  IV  NOT_4072(g4769,g3586);
  IV  NOT_4073(g5987,I9605);
  IV  NOT_4074(I11692,g7048);
  IV  NOT_4075(g7387,I11770);
  IV  NOT_4076(g11467,I17438);
  IV  NOT_4077(I9995,g5536);
  IV  NOT_4078(I12832,g7681);
  IV  NOT_4079(I4859,g578);
  IV  NOT_4080(I10051,g5702);
  IV  NOT_4081(I10072,g5719);
  IV  NOT_4082(g4212,I7453);
  IV  NOT_4083(I9479,g4954);
  IV  NOT_4084(g6689,g5830);
  IV  NOT_4085(g10130,I15392);
  IV  NOT_4086(g7756,I12433);
  IV  NOT_4087(g2297,g865);
  IV  NOT_4088(g11623,I17687);
  IV  NOT_4089(g6388,I10286);
  IV  NOT_4090(g10193,g10057);
  IV  NOT_4091(I16616,g10796);
  IV  NOT_4092(g11037,I16772);
  IV  NOT_4093(I10592,g5865);
  IV  NOT_4094(g5299,g4393);
  IV  NOT_4095(I10756,g5810);
  IV  NOT_4096(I15782,g10259);
  IV  NOT_4097(g7622,g7067);
  IV  NOT_4098(g3735,I6921);
  IV  NOT_4099(g7027,I11176);
  IV  NOT_4100(g7427,I11817);
  IV  NOT_4101(I17182,g11309);
  IV  NOT_4102(g10165,I15491);
  IV  NOT_4103(I13400,g8236);
  IV  NOT_4104(g10523,g10456);
  IV  NOT_4105(I17672,g11605);
  IV  NOT_4106(g3782,I7006);
  IV  NOT_4107(I13013,g8048);
  IV  NOT_4108(g5892,I9519);
  IV  NOT_4109(I11214,g6528);
  IV  NOT_4110(g7904,I12690);
  IV  NOT_4111(g11419,I17312);
  IV  NOT_4112(g2745,I5809);
  IV  NOT_4113(g2639,I5754);
  IV  NOT_4114(g6030,I9639);
  IV  NOT_4115(g2338,g1909);
  IV  NOT_4116(g11352,I17173);
  IV  NOT_4117(I15418,g10083);
  IV  NOT_4118(I5073,g34);
  IV  NOT_4119(I13329,g8116);
  IV  NOT_4120(I11207,g6524);
  IV  NOT_4121(g7446,g7148);
  IV  NOT_4122(g3475,g3056);
  IV  NOT_4123(I6999,g2905);
  IV  NOT_4124(g11155,g10950);
  IV  NOT_4125(I7284,g3255);
  IV  NOT_4126(I15266,g10001);
  IV  NOT_4127(g8990,I14391);
  IV  NOT_4128(I9156,g5032);
  IV  NOT_4129(I12099,g7258);
  IV  NOT_4130(I11005,g6386);
  IV  NOT_4131(I12388,g7219);
  IV  NOT_4132(I17331,g11357);
  IV  NOT_4133(I13005,g8046);
  IV  NOT_4134(g8888,I14232);
  IV  NOT_4135(g7403,I11783);
  IV  NOT_4136(g3627,I6784);
  IV  NOT_4137(g4822,g3706);
  IV  NOT_4138(g8029,I12871);
  IV  NOT_4139(g6564,g5784);
  IV  NOT_4140(I16808,g10906);
  IV  NOT_4141(g8171,I13068);
  IV  NOT_4142(g7345,I11683);
  IV  NOT_4143(I17513,g11482);
  IV  NOT_4144(I8711,g4530);
  IV  NOT_4145(g2808,g2156);
  IV  NOT_4146(g3292,g2373);
  IV  NOT_4147(I10846,g6729);
  IV  NOT_4148(g8787,I14094);
  IV  NOT_4149(I12251,g7076);
  IV  NOT_4150(g7763,I12454);
  IV  NOT_4151(I16101,g10381);
  IV  NOT_4152(g8956,I14319);
  IV  NOT_4153(g2707,g2041);
  IV  NOT_4154(I8827,g4477);
  IV  NOT_4155(g10437,g10333);
  IV  NOT_4156(I8133,g3632);
  IV  NOT_4157(g2759,I5843);
  IV  NOT_4158(I8333,g4456);
  IV  NOT_4159(I7420,g4167);
  IV  NOT_4160(g7637,I12251);
  IV  NOT_4161(I15589,g10161);
  IV  NOT_4162(g5078,g4372);
  IV  NOT_4163(g3039,g2310);
  IV  NOT_4164(g2201,g102);
  IV  NOT_4165(g3439,g3144);
  IV  NOT_4166(g7107,I11342);
  IV  NOT_4167(I7559,g4116);
  IV  NOT_4168(g7307,I11569);
  IV  NOT_4169(I12032,g6923);
  IV  NOT_4170(g8297,I13245);
  IV  NOT_4171(g10347,I15807);
  IV  NOT_4172(g5035,I8410);
  IV  NOT_4173(I6944,g2859);
  IV  NOT_4174(I8396,g4255);
  IV  NOT_4175(g10253,g10138);
  IV  NOT_4176(I6240,g878);
  IV  NOT_4177(I7931,g3624);
  IV  NOT_4178(g7359,I11725);
  IV  NOT_4179(g6108,I9779);
  IV  NOT_4180(g6308,I10183);
  IV  NOT_4181(I9810,g5576);
  IV  NOT_4182(g5082,g4840);
  IV  NOT_4183(g2449,g790);
  IV  NOT_4184(I9032,g4732);
  IV  NOT_4185(I11100,g6442);
  IV  NOT_4186(g5482,I8903);
  IV  NOT_4187(I14405,g8937);
  IV  NOT_4188(g10600,I16277);
  IV  NOT_4189(g11401,I17246);
  IV  NOT_4190(g10781,I16475);
  IV  NOT_4191(I4783,g873);
  IV  NOT_4192(I6043,g2267);
  IV  NOT_4193(I9053,g4752);
  IV  NOT_4194(g8684,I13969);
  IV  NOT_4195(g3583,I6742);
  IV  NOT_4196(g4895,I8250);
  IV  NOT_4197(g5876,g5361);
  IV  NOT_4198(g8138,I13013);
  IV  NOT_4199(I6443,g2363);
  IV  NOT_4200(I11235,g6538);
  IV  NOT_4201(g8338,I13394);
  IV  NOT_4202(g10236,g10190);
  IV  NOT_4203(g7757,I12436);
  IV  NOT_4204(g2604,I5713);
  IV  NOT_4205(g4062,I7185);
  IV  NOT_4206(g2098,I4938);
  IV  NOT_4207(I11683,g7069);
  IV  NOT_4208(g5656,I9129);
  IV  NOT_4209(g7416,I11800);
  IV  NOT_4210(g4620,I8031);
  IV  NOT_4211(g10351,I15817);
  IV  NOT_4212(g4462,I7825);
  IV  NOT_4213(I15864,g10339);
  IV  NOT_4214(I5399,g895);
  IV  NOT_4215(g6589,I10549);
  IV  NOT_4216(I12871,g7638);
  IV  NOT_4217(g10175,I15517);
  IV  NOT_4218(g10821,I16531);
  IV  NOT_4219(I7630,g3524);
  IV  NOT_4220(I15749,g10263);
  IV  NOT_4221(g2833,I5949);
  IV  NOT_4222(I6034,g2210);
  IV  NOT_4223(g7522,I11904);
  IV  NOT_4224(I8418,g4794);
  IV  NOT_4225(g7811,I12598);
  IV  NOT_4226(g7315,I11593);
  IV  NOT_4227(g11616,I17666);
  IV  NOT_4228(I17149,g11306);
  IV  NOT_4229(I6565,g2614);
  IV  NOT_4230(g7047,I11222);
  IV  NOT_4231(I7300,g2883);
  IV  NOT_4232(g11313,I17104);
  IV  NOT_4233(I12360,g7183);
  IV  NOT_4234(I8290,g4778);
  IV  NOT_4235(g10063,I15287);
  IV  NOT_4236(I17387,g11438);
  IV  NOT_4237(g8707,g8671);
  IV  NOT_4238(g6165,g5446);
  IV  NOT_4239(g10264,g10128);
  IV  NOT_4240(g6571,I10503);
  IV  NOT_4241(g6365,I10274);
  IV  NOT_4242(g6861,I10941);
  IV  NOT_4243(g5214,g4640);
  IV  NOT_4244(g10137,I15409);
  IV  NOT_4245(g6048,I9673);
  IV  NOT_4246(I11515,g6589);
  IV  NOT_4247(g9772,g9432);
  IV  NOT_4248(I11882,g6895);
  IV  NOT_4249(I5510,g588);
  IV  NOT_4250(g2539,I5652);
  IV  NOT_4251(g2896,g2356);
  IV  NOT_4252(I6347,g2462);
  IV  NOT_4253(I15704,g10238);
  IV  NOT_4254(I5245,g925);
  IV  NOT_4255(g6448,I10374);
  IV  NOT_4256(g9531,I14678);
  IV  NOT_4257(I15305,g10001);
  IV  NOT_4258(g6711,g5949);
  IV  NOT_4259(g6055,I9688);
  IV  NOT_4260(I12162,g7146);
  IV  NOT_4261(I17104,g11223);
  IV  NOT_4262(g10873,I16589);
  IV  NOT_4263(g11053,g10950);
  IV  NOT_4264(I8256,g4711);
  IV  NOT_4265(g9890,I15075);
  IV  NOT_4266(I10282,g6163);
  IV  NOT_4267(g3404,g3121);
  IV  NOT_4268(g6133,I9836);
  IV  NOT_4269(g11466,I17435);
  IV  NOT_4270(g5663,I9150);
  IV  NOT_4271(I10302,g6179);
  IV  NOT_4272(I6914,g2828);
  IV  NOT_4273(g9505,g9052);
  IV  NOT_4274(g2162,I5089);
  IV  NOT_4275(I7973,g3437);
  IV  NOT_4276(I15036,g9721);
  IV  NOT_4277(g2268,g654);
  IV  NOT_4278(g8449,I13645);
  IV  NOT_4279(g4192,I7393);
  IV  NOT_4280(I10105,g5736);
  IV  NOT_4281(g4298,g4130);
  IV  NOT_4282(g3764,I6971);
  IV  NOT_4283(I12451,g7538);
  IV  NOT_4284(g6846,I10910);
  IV  NOT_4285(g11036,I16769);
  IV  NOT_4286(I12472,g7539);
  IV  NOT_4287(g8575,I13816);
  IV  NOT_4288(g3546,g3307);
  IV  NOT_4289(I14105,g8776);
  IV  NOT_4290(g4485,g3546);
  IV  NOT_4291(I6013,g2200);
  IV  NOT_4292(g5402,I8842);
  IV  NOT_4293(g6196,g5446);
  IV  NOT_4294(g7880,g7479);
  IV  NOT_4295(g6396,I10296);
  IV  NOT_4296(g7595,I12123);
  IV  NOT_4297(g6803,I10819);
  IV  NOT_4298(g7537,I11947);
  IV  NOT_4299(g5236,g4361);
  IV  NOT_4300(I17368,g11423);
  IV  NOT_4301(g8604,g8479);
  IV  NOT_4302(g10208,I15580);
  IV  NOT_4303(I16239,g10525);
  IV  NOT_4304(g11642,I17730);
  IV  NOT_4305(g8498,g8353);
  IV  NOT_4306(I11584,g6827);
  IV  NOT_4307(g1972,g461);
  IV  NOT_4308(I8421,g4309);
  IV  NOT_4309(g9474,g9331);
  IV  NOT_4310(g7272,I11519);
  IV  NOT_4311(I13206,g8197);
  IV  NOT_4312(g10542,I16193);
  IV  NOT_4313(g6509,I10427);
  IV  NOT_4314(g11064,g10974);
  IV  NOT_4315(I15733,g10257);
  IV  NOT_4316(g7612,I12186);
  IV  NOT_4317(g7243,I11483);
  IV  NOT_4318(g2086,I4906);
  IV  NOT_4319(I11759,g7244);
  IV  NOT_4320(I11725,g7040);
  IV  NOT_4321(I12776,g7586);
  IV  NOT_4322(g5657,I9132);
  IV  NOT_4323(g10913,I16691);
  IV  NOT_4324(I16941,g11076);
  IV  NOT_4325(g2728,g2025);
  IV  NOT_4326(I13114,g7930);
  IV  NOT_4327(g6418,g6137);
  IV  NOT_4328(I11082,g6749);
  IV  NOT_4329(g7982,I12790);
  IV  NOT_4330(g4520,I7923);
  IV  NOT_4331(g5222,g4640);
  IV  NOT_4332(I17228,g11300);
  IV  NOT_4333(g11630,I17704);
  IV  NOT_4334(g2185,g46);
  IV  NOT_4335(g4219,g3635);
  IV  NOT_4336(g6290,I10129);
  IV  NOT_4337(I7151,g2642);
  IV  NOT_4338(g2881,I6031);
  IV  NOT_4339(I7351,g4061);
  IV  NOT_4340(I16518,g10718);
  IV  NOT_4341(I6601,g3186);
  IV  NOT_4342(I7648,g3727);
  IV  NOT_4343(I12825,g7696);
  IV  NOT_4344(g10320,I15756);
  IV  NOT_4345(g10905,I16667);
  IV  NOT_4346(g7629,I12229);
  IV  NOT_4347(I15665,g10193);
  IV  NOT_4348(g7328,I11632);
  IV  NOT_4349(g2070,g213);
  IV  NOT_4350(g10530,g10466);
  IV  NOT_4351(g3906,g3015);
  IV  NOT_4352(I17716,g11622);
  IV  NOT_4353(g7330,I11638);
  IV  NOT_4354(g10593,I16264);
  IV  NOT_4355(I4866,g579);
  IV  NOT_4356(g8362,I13466);
  IV  NOT_4357(I13744,g8297);
  IV  NOT_4358(g2025,g1696);
  IV  NOT_4359(I11345,g6692);
  IV  NOT_4360(g10346,I15804);
  IV  NOT_4361(I8631,g4425);
  IV  NOT_4362(g5899,g5361);
  IV  NOT_4363(g8419,I13571);
  IV  NOT_4364(g4958,I8328);
  IV  NOT_4365(g6256,I10027);
  IV  NOT_4366(g4176,I7345);
  IV  NOT_4367(g6816,I10858);
  IV  NOT_4368(g10122,I15374);
  IV  NOT_4369(g4376,I7691);
  IV  NOT_4370(g4005,I7143);
  IV  NOT_4371(g10464,I15983);
  IV  NOT_4372(I10027,g5751);
  IV  NOT_4373(I15476,g10114);
  IV  NOT_4374(I15485,g10092);
  IV  NOT_4375(g7800,I12565);
  IV  NOT_4376(g10034,I15238);
  IV  NOT_4377(g6181,g5426);
  IV  NOT_4378(I11804,g7190);
  IV  NOT_4379(I14249,g8804);
  IV  NOT_4380(g11454,I17419);
  IV  NOT_4381(g6847,g6482);
  IV  NOT_4382(g10292,I15698);
  IV  NOT_4383(I9475,g5445);
  IV  NOT_4384(I10248,g6125);
  IV  NOT_4385(g6685,I10648);
  IV  NOT_4386(g6197,I9930);
  IV  NOT_4387(g6700,g5949);
  IV  NOT_4388(I17112,g11227);
  IV  NOT_4389(I10710,g6088);
  IV  NOT_4390(g6397,I10299);
  IV  NOT_4391(I10003,g4908);
  IV  NOT_4392(g7213,I11447);
  IV  NOT_4393(I10204,g6031);
  IV  NOT_4394(I14552,g9264);
  IV  NOT_4395(I5336,g1700);
  IV  NOT_4396(g2131,I5060);
  IV  NOT_4397(g8486,g8348);
  IV  NOT_4398(I6784,g2742);
  IV  NOT_4399(g2006,g932);
  IV  NOT_4400(g2331,g658);
  IV  NOT_4401(I16577,g10825);
  IV  NOT_4402(g4733,I8089);
  IV  NOT_4403(g2406,g1365);
  IV  NOT_4404(g5844,I9461);
  IV  NOT_4405(I13332,g8206);
  IV  NOT_4406(g6263,I10048);
  IV  NOT_4407(g4270,g4013);
  IV  NOT_4408(I11135,g6679);
  IV  NOT_4409(I7372,g4057);
  IV  NOT_4410(g10136,I15406);
  IV  NOT_4411(g2635,g2003);
  IV  NOT_4412(I16439,g10702);
  IV  NOT_4413(I17742,g11636);
  IV  NOT_4414(I12318,g6862);
  IV  NOT_4415(g11074,g10901);
  IV  NOT_4416(g6950,I11094);
  IV  NOT_4417(g11239,g11112);
  IV  NOT_4418(I10081,g5735);
  IV  NOT_4419(I17096,g11219);
  IV  NOT_4420(g4225,I7478);
  IV  NOT_4421(I15238,g9974);
  IV  NOT_4422(g2087,g225);
  IV  NOT_4423(g11594,I17636);
  IV  NOT_4424(g3945,I7096);
  IV  NOT_4425(I7143,g2614);
  IV  NOT_4426(I5943,g2233);
  IV  NOT_4427(g2801,g2117);
  IV  NOT_4428(g5089,g4840);
  IV  NOT_4429(I13406,g8179);
  IV  NOT_4430(I9084,g4886);
  IV  NOT_4431(g3738,g3062);
  IV  NOT_4432(I13962,g8451);
  IV  NOT_4433(I14786,g9266);
  IV  NOT_4434(g7512,g7148);
  IV  NOT_4435(g8025,I12867);
  IV  NOT_4436(g9760,g9454);
  IV  NOT_4437(I6294,g2238);
  IV  NOT_4438(I17681,g11608);
  IV  NOT_4439(g8425,I13589);
  IV  NOT_4440(g3709,I6870);
  IV  NOT_4441(g4124,I7269);
  IV  NOT_4442(g4324,g4144);
  IV  NOT_4443(g2748,I5812);
  IV  NOT_4444(g6562,g5774);
  IV  NOT_4445(g7366,I11746);
  IV  NOT_4446(g10164,I15488);
  IV  NOT_4447(I11833,g7077);
  IV  NOT_4448(I11049,g6635);
  IV  NOT_4449(I15675,g10133);
  IV  NOT_4450(g4469,I7840);
  IV  NOT_4451(g5705,I9248);
  IV  NOT_4452(g5471,g4370);
  IV  NOT_4453(g2755,I5833);
  IV  NOT_4454(g11185,I16956);
  IV  NOT_4455(g7056,I11249);
  IV  NOT_4456(I17730,g11638);
  IV  NOT_4457(g3907,I7076);
  IV  NOT_4458(g10891,I16635);
  IV  NOT_4459(g2226,g86);
  IV  NOT_4460(I6501,g2578);
  IV  NOT_4461(I10090,g5767);
  IV  NOT_4462(g6723,I10716);
  IV  NOT_4463(I13048,g8059);
  IV  NOT_4464(g6257,I10030);
  IV  NOT_4465(I14090,g8771);
  IV  NOT_4466(g11518,I17563);
  IV  NOT_4467(g4177,I7348);
  IV  NOT_4468(I6156,g2119);
  IV  NOT_4469(g6101,I9762);
  IV  NOT_4470(g7148,I11397);
  IV  NOT_4471(g6817,I10861);
  IV  NOT_4472(g7649,I12258);
  IV  NOT_4473(g5948,I9588);
  IV  NOT_4474(g6301,I10162);
  IV  NOT_4475(g7348,I11692);
  IV  NOT_4476(I6356,g2459);
  IV  NOT_4477(g4377,I7694);
  IV  NOT_4478(g4206,I7435);
  IV  NOT_4479(I10651,g6035);
  IV  NOT_4480(g3517,I6702);
  IV  NOT_4481(g10575,g10523);
  IV  NOT_4482(I14182,g8788);
  IV  NOT_4483(I14672,g9261);
  IV  NOT_4484(g7355,I11713);
  IV  NOT_4485(g2045,g1811);
  IV  NOT_4486(g7851,g7479);
  IV  NOT_4487(I17549,g11501);
  IV  NOT_4488(g3876,I7061);
  IV  NOT_4489(g8131,g8020);
  IV  NOT_4490(g10327,I15771);
  IV  NOT_4491(g8331,I13373);
  IV  NOT_4492(g2173,I5120);
  IV  NOT_4493(I12120,g7106);
  IV  NOT_4494(g2373,g471);
  IV  NOT_4495(g4287,I7546);
  IV  NOT_4496(I9276,g5241);
  IV  NOT_4497(g10537,I16178);
  IV  NOT_4498(I10331,g6198);
  IV  NOT_4499(g7964,g7651);
  IV  NOT_4500(g8635,I13918);
  IV  NOT_4501(g6751,I10762);
  IV  NOT_4502(I12562,g7377);
  IV  NOT_4503(I8011,g3820);
  IV  NOT_4504(I11947,g6905);
  IV  NOT_4505(g8105,g7992);
  IV  NOT_4506(g2169,g42);
  IV  NOT_4507(I5395,g892);
  IV  NOT_4508(I14449,g8973);
  IV  NOT_4509(g10283,g10166);
  IV  NOT_4510(g2369,g617);
  IV  NOT_4511(I5913,g2169);
  IV  NOT_4512(I11106,g6667);
  IV  NOT_4513(g8487,g8350);
  IV  NOT_4514(g2602,I5707);
  IV  NOT_4515(I11605,g6834);
  IV  NOT_4516(g4199,I7414);
  IV  NOT_4517(g6585,I10541);
  IV  NOT_4518(g2007,g936);
  IV  NOT_4519(g5773,I9359);
  IV  NOT_4520(g10492,I16111);
  IV  NOT_4521(g4399,g3638);
  IV  NOT_4522(g7463,g6921);
  IV  NOT_4523(g2407,g197);
  IV  NOT_4524(I6163,g2547);
  IV  NOT_4525(g2920,g2462);
  IV  NOT_4526(I14961,g9769);
  IV  NOT_4527(g2578,g1962);
  IV  NOT_4528(g2868,I6010);
  IV  NOT_4529(g3214,I6391);
  IV  NOT_4530(g4781,I8147);
  IV  NOT_4531(g6041,I9658);
  IV  NOT_4532(I6363,g2459);
  IV  NOT_4533(I7202,g2647);
  IV  NOT_4534(I15729,g10254);
  IV  NOT_4535(I13812,g8519);
  IV  NOT_4536(I9647,g5148);
  IV  NOT_4537(g4898,I8259);
  IV  NOT_4538(g6441,g6151);
  IV  NOT_4539(I13463,g8156);
  IV  NOT_4540(g9451,I14642);
  IV  NOT_4541(g4900,I8265);
  IV  NOT_4542(I6432,g2350);
  IV  NOT_4543(g11501,I17522);
  IV  NOT_4544(g3110,g2482);
  IV  NOT_4545(g11577,I17613);
  IV  NOT_4546(g7279,g6382);
  IV  NOT_4547(g5836,g5320);
  IV  NOT_4548(g4510,I7909);
  IV  NOT_4549(g11439,I17368);
  IV  NOT_4550(g3663,I6832);
  IV  NOT_4551(I12427,g7636);
  IV  NOT_4552(g10091,I15320);
  IV  NOT_4553(g9346,I14543);
  IV  NOT_4554(I12366,g7134);
  IV  NOT_4555(g2261,g1713);
  IV  NOT_4556(g7619,I12205);
  IV  NOT_4557(g7318,I11602);
  IV  NOT_4558(g2793,g2276);
  IV  NOT_4559(g4291,g4013);
  IV  NOT_4560(g7872,I12655);
  IV  NOT_4561(g11438,I17365);
  IV  NOT_4562(g10174,I15514);
  IV  NOT_4563(g10796,I16500);
  IV  NOT_4564(I16664,g10795);
  IV  NOT_4565(g9103,g8892);
  IV  NOT_4566(I8080,g3538);
  IV  NOT_4567(g2015,g1107);
  IV  NOT_4568(g6368,g5987);
  IV  NOT_4569(g8445,I13633);
  IV  NOT_4570(I7776,g3773);
  IV  NOT_4571(g7057,I11252);
  IV  NOT_4572(g2227,g95);
  IV  NOT_4573(g4344,g3946);
  IV  NOT_4574(I5142,g639);
  IV  NOT_4575(I7593,g4142);
  IV  NOT_4576(I5248,g1110);
  IV  NOT_4577(g7989,I12805);
  IV  NOT_4578(I9224,g5063);
  IV  NOT_4579(I15284,g10034);
  IV  NOT_4580(g3762,I6965);
  IV  NOT_4581(I12403,g7611);
  IV  NOT_4582(I12547,g7673);
  IV  NOT_4583(g4207,I7438);
  IV  NOT_4584(g11083,g10913);
  IV  NOT_4585(g11348,g11276);
  IV  NOT_4586(g10390,g10309);
  IV  NOT_4587(I16484,g10770);
  IV  NOT_4588(g9732,I14873);
  IV  NOT_4589(I5815,g1994);
  IV  NOT_4590(I9120,g5218);
  IV  NOT_4591(g11284,g11208);
  IV  NOT_4592(I9320,g5013);
  IV  NOT_4593(g2246,g1810);
  IV  NOT_4594(g5822,g5320);
  IV  NOT_4595(g4819,g3354);
  IV  NOT_4596(g3877,I7064);
  IV  NOT_4597(g9508,g9271);
  IV  NOT_4598(I12226,g7066);
  IV  NOT_4599(g8007,I12843);
  IV  NOT_4600(I7264,g3252);
  IV  NOT_4601(g11622,I17684);
  IV  NOT_4602(g2203,g677);
  IV  NOT_4603(g7686,g7148);
  IV  NOT_4604(g10192,I15554);
  IV  NOT_4605(I10620,g5884);
  IV  NOT_4606(I5497,g587);
  IV  NOT_4607(I6929,g2846);
  IV  NOT_4608(I12481,g7570);
  IV  NOT_4609(I13421,g8200);
  IV  NOT_4610(I16200,g10494);
  IV  NOT_4611(g8868,I14176);
  IV  NOT_4612(I5960,g2239);
  IV  NOT_4613(I7360,g4081);
  IV  NOT_4614(I14097,g8773);
  IV  NOT_4615(I9617,g5405);
  IV  NOT_4616(g6856,I10924);
  IV  NOT_4617(g6411,g6135);
  IV  NOT_4618(g6734,I10733);
  IV  NOT_4619(I9789,g5401);
  IV  NOT_4620(I10343,g6003);
  IV  NOT_4621(g8535,I13744);
  IV  NOT_4622(I7450,g3704);
  IV  NOT_4623(I10971,g6344);
  IV  NOT_4624(g7321,I11611);
  IV  NOT_4625(g8582,I13825);
  IV  NOT_4626(g7670,I12289);
  IV  NOT_4627(I17261,g11346);
  IV  NOT_4628(g4215,I7462);
  IV  NOT_4629(I7996,g3462);
  IV  NOT_4630(g11653,I17761);
  IV  NOT_4631(g2502,I5579);
  IV  NOT_4632(g4886,I8231);
  IV  NOT_4633(g4951,I8320);
  IV  NOT_4634(I16799,g11017);
  IV  NOT_4635(g7232,I11472);
  IV  NOT_4636(I12490,g7637);
  IV  NOT_4637(g10553,I16220);
  IV  NOT_4638(g8015,I12857);
  IV  NOT_4639(I15415,g10075);
  IV  NOT_4640(g5895,g5361);
  IV  NOT_4641(g7938,g7403);
  IV  NOT_4642(I8126,g3662);
  IV  NOT_4643(g7813,I12604);
  IV  NOT_4644(I5979,g2543);
  IV  NOT_4645(g4314,g4013);
  IV  NOT_4646(I5218,g1104);
  IV  NOT_4647(g5062,g4840);
  IV  NOT_4648(I13788,g8517);
  IV  NOT_4649(g9347,I14546);
  IV  NOT_4650(I12376,g7195);
  IV  NOT_4651(g10326,I15768);
  IV  NOT_4652(g5620,g4417);
  IV  NOT_4653(g7909,g7664);
  IV  NOT_4654(g2689,g2038);
  IV  NOT_4655(I12103,g6859);
  IV  NOT_4656(I11829,g7213);
  IV  NOT_4657(g6863,g6740);
  IV  NOT_4658(I16184,g10484);
  IV  NOT_4659(I16805,g10904);
  IV  NOT_4660(g10536,I16175);
  IV  NOT_4661(g8664,I13949);
  IV  NOT_4662(g10040,I15247);
  IV  NOT_4663(I10412,g5821);
  IV  NOT_4664(I12354,g7143);
  IV  NOT_4665(g2216,g41);
  IV  NOT_4666(g9533,I14684);
  IV  NOT_4667(g6713,I10698);
  IV  NOT_4668(I14412,g8939);
  IV  NOT_4669(g7519,g6956);
  IV  NOT_4670(I13828,g8488);
  IV  NOT_4671(g10904,I16664);
  IV  NOT_4672(g2028,g1703);
  IV  NOT_4673(I14133,g8772);
  IV  NOT_4674(g10252,g10137);
  IV  NOT_4675(g8721,g8582);
  IV  NOT_4676(g6569,I10499);
  IV  NOT_4677(g10621,I16298);
  IV  NOT_4678(g7606,I12168);
  IV  NOT_4679(I6894,g2813);
  IV  NOT_4680(I13344,g8121);
  IV  NOT_4681(I10228,g6113);
  IV  NOT_4682(g2247,I5258);
  IV  NOT_4683(I14228,g8797);
  IV  NOT_4684(g4336,g4130);
  IV  NOT_4685(g3394,I6598);
  IV  NOT_4686(I5830,g2067);
  IV  NOT_4687(g2564,g1814);
  IV  NOT_4688(g7687,I12318);
  IV  NOT_4689(g4768,I8126);
  IV  NOT_4690(g11576,I17610);
  IV  NOT_4691(I10716,g6093);
  IV  NOT_4692(I13682,g8310);
  IV  NOT_4693(g3731,I6911);
  IV  NOT_4694(I15554,g10088);
  IV  NOT_4695(g2826,g2163);
  IV  NOT_4696(I6661,g2752);
  IV  NOT_4697(g6688,I10655);
  IV  NOT_4698(I11173,g6500);
  IV  NOT_4699(g10183,g10042);
  IV  NOT_4700(g6857,I10927);
  IV  NOT_4701(g5192,g4640);
  IV  NOT_4702(g5085,g4377);
  IV  NOT_4703(I5221,g1407);
  IV  NOT_4704(g9820,I14961);
  IV  NOT_4705(g4943,I8311);
  IV  NOT_4706(I12190,g7268);
  IV  NOT_4707(I7674,g3352);
  IV  NOT_4708(g11200,g11112);
  IV  NOT_4709(g10062,I15284);
  IV  NOT_4710(g3705,g3113);
  IV  NOT_4711(I16214,g10500);
  IV  NOT_4712(I17271,g11388);
  IV  NOT_4713(I12520,g7415);
  IV  NOT_4714(g2638,I5751);
  IV  NOT_4715(g4065,g2794);
  IV  NOT_4716(I8161,g3637);
  IV  NOT_4717(g4887,I8234);
  IV  NOT_4718(g4228,g3914);
  IV  NOT_4719(g4322,I7593);
  IV  NOT_4720(g7570,I12032);
  IV  NOT_4721(g2108,I4992);
  IV  NOT_4722(g5941,I9571);
  IV  NOT_4723(I14379,g8961);
  IV  NOT_4724(g2609,I5728);
  IV  NOT_4725(g4934,g4243);
  IV  NOT_4726(g7341,I11671);
  IV  NOT_4727(I11029,g6485);
  IV  NOT_4728(g10851,I16553);
  IV  NOT_4729(g10872,I16586);
  IV  NOT_4730(g11052,I16817);
  IV  NOT_4731(I5932,g2539);
  IV  NOT_4732(I10958,g6559);
  IV  NOT_4733(g6400,I10308);
  IV  NOT_4734(I14112,g8777);
  IV  NOT_4735(I10378,g6244);
  IV  NOT_4736(g7525,I11921);
  IV  NOT_4737(I7680,g3736);
  IV  NOT_4738(I14958,g9767);
  IV  NOT_4739(g2883,I6037);
  IV  NOT_4740(g8671,I13956);
  IV  NOT_4741(I6484,g2073);
  IV  NOT_4742(I6439,g2352);
  IV  NOT_4743(I9915,g5304);
  IV  NOT_4744(g3254,g2322);
  IV  NOT_4745(g9775,g9474);
  IV  NOT_4746(I17736,g11640);
  IV  NOT_4747(I15798,g10281);
  IV  NOT_4748(g3814,g3228);
  IV  NOT_4749(g5708,I9253);
  IV  NOT_4750(I10096,g5794);
  IV  NOT_4751(g2217,I5192);
  IV  NOT_4752(g2758,I5840);
  IV  NOT_4753(g5520,I8943);
  IV  NOT_4754(I14944,g9454);
  IV  NOT_4755(I17198,g11319);
  IV  NOT_4756(I15184,g9974);
  IV  NOT_4757(g4096,I7236);
  IV  NOT_4758(g8564,I13785);
  IV  NOT_4759(g3038,g1982);
  IV  NOT_4760(g4496,I7889);
  IV  NOT_4761(I8303,g4784);
  IV  NOT_4762(g11184,I16953);
  IV  NOT_4763(g5252,g4640);
  IV  NOT_4764(g7607,I12171);
  IV  NOT_4765(I17528,g11487);
  IV  NOT_4766(I6702,g2801);
  IV  NOT_4767(g3773,I6996);
  IV  NOT_4768(g5812,g5320);
  IV  NOT_4769(g3009,g2135);
  IV  NOT_4770(I14681,g9110);
  IV  NOT_4771(g2165,I5098);
  IV  NOT_4772(g6183,g5320);
  IV  NOT_4773(g2571,g1822);
  IV  NOT_4774(g7659,I12274);
  IV  NOT_4775(g2861,I6001);
  IV  NOT_4776(g7358,I11722);
  IV  NOT_4777(g4195,I7402);
  IV  NOT_4778(g5176,g4682);
  IV  NOT_4779(g6220,g5446);
  IV  NOT_4780(I5716,g2068);
  IV  NOT_4781(g10574,I16239);
  IV  NOT_4782(I17764,g11651);
  IV  NOT_4783(I5149,g1453);
  IV  NOT_4784(g4395,I7732);
  IV  NOT_4785(g10047,I15266);
  IV  NOT_4786(g4337,g4144);
  IV  NOT_4787(g4913,I8285);
  IV  NOT_4788(I17365,g11380);
  IV  NOT_4789(I14802,g9666);
  IV  NOT_4790(g10205,g10176);
  IV  NOT_4791(g2055,g1950);
  IV  NOT_4792(g3769,I6982);
  IV  NOT_4793(g10912,I16688);
  IV  NOT_4794(g10311,g10242);
  IV  NOT_4795(g2455,g826);
  IV  NOT_4796(g9739,I14884);
  IV  NOT_4797(g2827,g2164);
  IV  NOT_4798(I6952,g2867);
  IV  NOT_4799(I14793,g9269);
  IV  NOT_4800(g3212,I6385);
  IV  NOT_4801(I9402,g5107);
  IV  NOT_4802(I12339,g7054);
  IV  NOT_4803(I8240,g4380);
  IV  NOT_4804(g1975,g622);
  IV  NOT_4805(I5198,g143);
  IV  NOT_4806(I12296,g7236);
  IV  NOT_4807(g7311,I11581);
  IV  NOT_4808(g2774,g2276);
  IV  NOT_4809(I6616,g3186);
  IV  NOT_4810(g3967,g3247);
  IV  NOT_4811(I17161,g11314);
  IV  NOT_4812(g6588,I10546);
  IV  NOT_4813(I4935,g585);
  IV  NOT_4814(I12644,g7729);
  IV  NOT_4815(g2846,I5970);
  IV  NOT_4816(I9762,g5276);
  IV  NOT_4817(I10549,g6184);
  IV  NOT_4818(g9079,g8892);
  IV  NOT_4819(I13648,g8376);
  IV  NOT_4820(g10051,I15272);
  IV  NOT_4821(I14690,g9150);
  IV  NOT_4822(g6161,I9886);
  IV  NOT_4823(I14549,g9262);
  IV  NOT_4824(g7615,I12193);
  IV  NOT_4825(g6361,g5867);
  IV  NOT_4826(g2196,g91);
  IV  NOT_4827(g4266,g3688);
  IV  NOT_4828(I7600,g4159);
  IV  NOT_4829(g9668,g9490);
  IV  NOT_4830(g2396,g1389);
  IV  NOT_4831(g10592,I16261);
  IV  NOT_4832(I15400,g10069);
  IV  NOT_4833(g2803,g2154);
  IV  NOT_4834(g5733,I9287);
  IV  NOT_4835(I17225,g11298);
  IV  NOT_4836(g11400,I17243);
  IV  NOT_4837(g6051,I9680);
  IV  NOT_4838(I11770,g7202);
  IV  NOT_4839(g5270,g4367);
  IV  NOT_4840(g7374,I11752);
  IV  NOT_4841(I11563,g6819);
  IV  NOT_4842(I8116,g3627);
  IV  NOT_4843(g6127,I9826);
  IV  NOT_4844(g6451,I10381);
  IV  NOT_4845(g8758,I14055);
  IV  NOT_4846(g8066,I12916);
  IV  NOT_4847(g8589,I13834);
  IV  NOT_4848(I15329,g9995);
  IV  NOT_4849(g7985,I12799);
  IV  NOT_4850(I17258,g11345);
  IV  NOT_4851(g4142,I7288);
  IV  NOT_4852(g2509,I5588);
  IV  NOT_4853(I16407,g10696);
  IV  NOT_4854(I15539,g10069);
  IV  NOT_4855(I6546,g2987);
  IV  NOT_4856(g5073,g4840);
  IV  NOT_4857(g10350,I15814);
  IV  NOT_4858(g11207,I16982);
  IV  NOT_4859(g1984,g758);
  IV  NOT_4860(I10317,g6003);
  IV  NOT_4861(g7284,I11528);
  IV  NOT_4862(g11539,g11519);
  IV  NOT_4863(g6146,I9863);
  IV  NOT_4864(g10820,I16528);
  IV  NOT_4865(g4081,I7210);
  IV  NOT_4866(g7545,I11967);
  IV  NOT_4867(g9356,I14573);
  IV  NOT_4868(g8571,I13806);
  IV  NOT_4869(I8147,g3633);
  IV  NOT_4870(g2662,g2014);
  IV  NOT_4871(g5124,g4596);
  IV  NOT_4872(g2018,g1336);
  IV  NOT_4873(g5980,I9594);
  IV  NOT_4874(g2067,g108);
  IV  NOT_4875(g7380,g7279);
  IV  NOT_4876(g8448,I13642);
  IV  NOT_4877(g6103,I9766);
  IV  NOT_4878(I10129,g5688);
  IV  NOT_4879(I9930,g5317);
  IV  NOT_4880(I11767,g7201);
  IV  NOT_4881(I11794,g7188);
  IV  NOT_4882(g8711,g8677);
  IV  NOT_4883(g7591,I12103);
  IV  NOT_4884(g6303,I10168);
  IV  NOT_4885(g2418,I5497);
  IV  NOT_4886(I11845,g6869);
  IV  NOT_4887(g5069,g4368);
  IV  NOT_4888(I13794,g8472);
  IV  NOT_4889(I10057,g5741);
  IV  NOT_4890(g4726,g3546);
  IV  NOT_4891(g2994,g2057);
  IV  NOT_4892(g5469,I8880);
  IV  NOT_4893(g7853,I12652);
  IV  NOT_4894(g4354,I7639);
  IV  NOT_4895(I5258,g67);
  IV  NOT_4896(g7020,I11159);
  IV  NOT_4897(I5818,g2098);
  IV  NOT_4898(g8133,I13002);
  IV  NOT_4899(g8333,I13379);
  IV  NOT_4900(g7420,I11804);
  IV  NOT_4901(I15241,g10013);
  IV  NOT_4902(I11898,g6896);
  IV  NOT_4903(g5177,g4596);
  IV  NOT_4904(g6732,I10729);
  IV  NOT_4905(I12867,g7638);
  IV  NOT_4906(I17657,g11598);
  IV  NOT_4907(I13633,g8346);
  IV  NOT_4908(g11241,g11112);
  IV  NOT_4909(I16206,g10453);
  IV  NOT_4910(I10299,g6243);
  IV  NOT_4911(g2256,I5279);
  IV  NOT_4912(I11191,g6514);
  IV  NOT_4913(I11719,g7029);
  IV  NOT_4914(g7559,I12009);
  IV  NOT_4915(I14323,g8817);
  IV  NOT_4916(g10691,I16360);
  IV  NOT_4917(g7794,I12547);
  IV  NOT_4918(I7076,g2985);
  IV  NOT_4919(I13191,g8132);
  IV  NOT_4920(I14299,g8810);
  IV  NOT_4921(I7889,g3373);
  IV  NOT_4922(g8196,I13125);
  IV  NOT_4923(g6944,I11082);
  IV  NOT_4924(g8803,I14130);
  IV  NOT_4925(I6277,g1206);
  IV  NOT_4926(g6072,g4977);
  IV  NOT_4927(I15771,g10250);
  IV  NOT_4928(I9237,g5205);
  IV  NOT_4929(I17337,g11363);
  IV  NOT_4930(g2181,I5142);
  IV  NOT_4931(g8538,I13747);
  IV  NOT_4932(g2381,g1368);
  IV  NOT_4933(g9432,g9313);
  IV  NOT_4934(I15235,g9968);
  IV  NOT_4935(I6789,g2748);
  IV  NOT_4936(I16114,g10387);
  IV  NOT_4937(g4783,g3829);
  IV  NOT_4938(g6043,I9662);
  IV  NOT_4939(I12910,g7922);
  IV  NOT_4940(I7375,g4062);
  IV  NOT_4941(g2847,I5973);
  IV  NOT_4942(g8780,I14077);
  IV  NOT_4943(g6443,g6157);
  IV  NOT_4944(I12202,g6983);
  IV  NOT_4945(g8509,g8366);
  IV  NOT_4946(g9453,g9100);
  IV  NOT_4947(g4112,g2994);
  IV  NOT_4948(g7905,g7450);
  IV  NOT_4949(g2197,g101);
  IV  NOT_4950(I7651,g3332);
  IV  NOT_4951(g4312,g4144);
  IV  NOT_4952(I8820,g4473);
  IV  NOT_4953(I11440,g6577);
  IV  NOT_4954(g10929,g10827);
  IV  NOT_4955(I12496,g7724);
  IV  NOT_4956(g2021,g1341);
  IV  NOT_4957(I9194,g5236);
  IV  NOT_4958(g7628,I12226);
  IV  NOT_4959(I9394,g5195);
  IV  NOT_4960(g6116,I9801);
  IV  NOT_4961(g2421,g1374);
  IV  NOT_4962(g7630,I12232);
  IV  NOT_4963(g4001,g3200);
  IV  NOT_4964(I12978,g8040);
  IV  NOT_4965(I14232,g8800);
  IV  NOT_4966(g10928,g10827);
  IV  NOT_4967(g8067,I12919);
  IV  NOT_4968(I9731,g5255);
  IV  NOT_4969(g5898,g5361);
  IV  NOT_4970(g8418,I13568);
  IV  NOT_4971(g6434,I10352);
  IV  NOT_4972(g4676,g3354);
  IV  NOT_4973(g5900,I9531);
  IV  NOT_4974(g6565,g5790);
  IV  NOT_4975(I5821,g2101);
  IV  NOT_4976(I6299,g2242);
  IV  NOT_4977(I11926,g6900);
  IV  NOT_4978(g8290,I13224);
  IV  NOT_4979(I12986,g8042);
  IV  NOT_4980(g4129,I7280);
  IV  NOT_4981(g5797,I9399);
  IV  NOT_4982(g4329,g4144);
  IV  NOT_4983(I14697,g9260);
  IV  NOT_4984(g4761,g3440);
  IV  NOT_4985(g11515,g11490);
  IV  NOT_4986(I7384,g4082);
  IV  NOT_4987(I13612,g8325);
  IV  NOT_4988(g5245,g4369);
  IV  NOT_4989(I7339,g4004);
  IV  NOT_4990(I13099,g7927);
  IV  NOT_4991(I12384,g7212);
  IV  NOT_4992(g8093,I12948);
  IV  NOT_4993(I13388,g8230);
  IV  NOT_4994(g6681,g5830);
  IV  NOT_4995(I11701,g7065);
  IV  NOT_4996(I11534,g6917);
  IV  NOT_4997(g10787,I16487);
  IV  NOT_4998(g5291,g4384);
  IV  NOT_4999(g3392,g3121);
  IV  NOT_5000(I11272,g6546);
  IV  NOT_5001(g10282,g10164);
  IV  NOT_5002(g7750,I12415);
  IV  NOT_5003(g3485,g2662);
  IV  NOT_5004(g2562,g1383);
  IV  NOT_5005(g6697,g5949);
  IV  NOT_5006(g5144,g4682);
  IV  NOT_5007(g4592,g3829);
  IV  NOT_5008(g6914,I11024);
  IV  NOT_5009(I17444,g11446);
  IV  NOT_5010(g5344,I8811);
  IV  NOT_5011(g6210,g5205);
  IV  NOT_5012(I12150,g7074);
  IV  NOT_5013(g4746,I8098);
  IV  NOT_5014(g8181,I13096);
  IV  NOT_5015(g10827,I16543);
  IV  NOT_5016(g6596,I10566);
  IV  NOT_5017(I6738,g3113);
  IV  NOT_5018(g4221,g3914);
  IV  NOT_5019(g8381,I13489);
  IV  NOT_5020(g2101,I4951);
  IV  NOT_5021(g2817,I5919);
  IV  NOT_5022(g3941,g3015);
  IV  NOT_5023(g7040,I11207);
  IV  NOT_5024(g6413,I10325);
  IV  NOT_5025(I10831,g6710);
  IV  NOT_5026(g7440,I11836);
  IV  NOT_5027(g8197,I13128);
  IV  NOT_5028(g8700,g8574);
  IV  NOT_5029(I10445,g5770);
  IV  NOT_5030(I7523,g4095);
  IV  NOT_5031(I11140,g6448);
  IV  NOT_5032(I12196,g7272);
  IV  NOT_5033(g2605,I5716);
  IV  NOT_5034(g11441,I17374);
  IV  NOT_5035(I9150,g5012);
  IV  NOT_5036(I10499,g6149);
  IV  NOT_5037(g8421,I13577);
  IV  NOT_5038(g7123,I11360);
  IV  NOT_5039(g5088,I8456);
  IV  NOT_5040(g11206,I16979);
  IV  NOT_5041(g7323,I11617);
  IV  NOT_5042(I14499,g8889);
  IV  NOT_5043(I6907,g2994);
  IV  NOT_5044(I12526,g7648);
  IV  NOT_5045(g10803,g10708);
  IV  NOT_5046(I7205,g2632);
  IV  NOT_5047(I9773,g4934);
  IV  NOT_5048(I15759,g10267);
  IV  NOT_5049(I11061,g6641);
  IV  NOT_5050(I15725,g10251);
  IV  NOT_5051(g5701,I9240);
  IV  NOT_5052(g3708,I6867);
  IV  NOT_5053(g4953,I8324);
  IV  NOT_5054(g2751,I5821);
  IV  NOT_5055(g3520,g2779);
  IV  NOT_5056(g8950,I14303);
  IV  NOT_5057(I16500,g10711);
  IV  NOT_5058(g3219,I6395);
  IV  NOT_5059(I6517,g3271);
  IV  NOT_5060(I6690,g2743);
  IV  NOT_5061(I9409,g5013);
  IV  NOT_5062(I15114,g9875);
  IV  NOT_5063(I5427,g913);
  IV  NOT_5064(g4468,I7837);
  IV  NOT_5065(I15082,g9719);
  IV  NOT_5066(g6117,I9804);
  IV  NOT_5067(I14989,g9813);
  IV  NOT_5068(I17158,g11312);
  IV  NOT_5069(g3252,I6414);
  IV  NOT_5070(g10881,I16613);
  IV  NOT_5071(I7104,g3186);
  IV  NOT_5072(g11435,I17356);
  IV  NOT_5073(I6876,g2956);
  IV  NOT_5074(I9769,g5287);
  IV  NOT_5075(g11082,I16859);
  IV  NOT_5076(g3812,g3228);
  IV  NOT_5077(I7099,g3228);
  IV  NOT_5078(I12457,g7559);
  IV  NOT_5079(I10924,g6736);
  IV  NOT_5080(g5886,g5361);
  IV  NOT_5081(g11107,g10974);
  IV  NOT_5082(I9836,g5405);
  IV  NOT_5083(I14080,g8714);
  IV  NOT_5084(g7351,I11701);
  IV  NOT_5085(g2041,g1791);
  IV  NOT_5086(g7648,I12255);
  IV  NOT_5087(g7530,I11926);
  IV  NOT_5088(I11360,g6351);
  IV  NOT_5089(g8562,I13779);
  IV  NOT_5090(I15744,g10261);
  IV  NOT_5091(I13360,g8126);
  IV  NOT_5092(I17353,g11381);
  IV  NOT_5093(g3405,g3144);
  IV  NOT_5094(g5114,I8506);
  IV  NOT_5095(I5403,g636);
  IV  NOT_5096(g9778,g9474);
  IV  NOT_5097(g5314,g4387);
  IV  NOT_5098(I11447,g6431);
  IV  NOT_5099(g11345,I17158);
  IV  NOT_5100(g9894,I15085);
  IV  NOT_5101(g8723,g8585);
  IV  NOT_5102(g4716,g3546);
  IV  NOT_5103(I11162,g6479);
  IV  NOT_5104(I16613,g10794);
  IV  NOT_5105(g11399,I17240);
  IV  NOT_5106(g3765,g3120);
  IV  NOT_5107(I10753,g5814);
  IV  NOT_5108(I10461,g5849);
  IV  NOT_5109(I5391,g1101);
  IV  NOT_5110(g3911,g3015);
  IV  NOT_5111(I9229,g4954);
  IV  NOT_5112(g7010,I11155);
  IV  NOT_5113(g6581,I10531);
  IV  NOT_5114(g10890,I16632);
  IV  NOT_5115(g5650,I9111);
  IV  NOT_5116(g7410,I11790);
  IV  NOT_5117(g9782,I14933);
  IV  NOT_5118(g11398,I17237);
  IV  NOT_5119(I15804,g10283);
  IV  NOT_5120(I16947,g11080);
  IV  NOT_5121(I5695,g575);
  IV  NOT_5122(g10249,g10135);
  IV  NOT_5123(g2168,I5111);
  IV  NOT_5124(g2669,g2015);
  IV  NOT_5125(g6060,I9695);
  IV  NOT_5126(I16273,g10559);
  IV  NOT_5127(g2368,I5445);
  IV  NOT_5128(I11629,g6914);
  IV  NOT_5129(g11652,I17758);
  IV  NOT_5130(I9822,g5219);
  IV  NOT_5131(g9661,I14786);
  IV  NOT_5132(g4198,I7411);
  IV  NOT_5133(g4747,g3586);
  IV  NOT_5134(I11472,g6488);
  IV  NOT_5135(I10736,g6104);
  IV  NOT_5136(g4398,g3914);
  IV  NOT_5137(I13451,g8152);
  IV  NOT_5138(g3733,I6917);
  IV  NOT_5139(I7444,g3683);
  IV  NOT_5140(g10248,g10134);
  IV  NOT_5141(g2772,g2508);
  IV  NOT_5142(I7269,g2851);
  IV  NOT_5143(I15263,g9995);
  IV  NOT_5144(I10198,g6118);
  IV  NOT_5145(I12300,g7240);
  IV  NOT_5146(g10552,I16217);
  IV  NOT_5147(g8751,g8632);
  IV  NOT_5148(I15332,g10001);
  IV  NOT_5149(g10204,g10174);
  IV  NOT_5150(g2743,I5801);
  IV  NOT_5151(g4241,g3664);
  IV  NOT_5152(g2890,I6052);
  IV  NOT_5153(g5768,I9352);
  IV  NOT_5154(I10843,g6723);
  IV  NOT_5155(g8585,I13828);
  IV  NOT_5156(I5858,g2529);
  IV  NOT_5157(g5594,I9016);
  IV  NOT_5158(I14528,g9270);
  IV  NOT_5159(g3473,I6676);
  IV  NOT_5160(g7278,I11524);
  IV  NOT_5161(I14330,g8819);
  IV  NOT_5162(g9526,g9256);
  IV  NOT_5163(I4938,g261);
  IV  NOT_5164(I8250,g4589);
  IV  NOT_5165(I11071,g6656);
  IV  NOT_5166(I15406,g10065);
  IV  NOT_5167(I15962,g10405);
  IV  NOT_5168(g2011,g976);
  IV  NOT_5169(g6995,g6482);
  IV  NOT_5170(g7618,I12202);
  IV  NOT_5171(g3980,g3121);
  IV  NOT_5172(g8441,I13621);
  IV  NOT_5173(g11406,I17261);
  IV  NOT_5174(g5943,I9581);
  IV  NOT_5175(g7343,I11677);
  IV  NOT_5176(g2411,I5494);
  IV  NOT_5177(I10132,g5696);
  IV  NOT_5178(g10786,I16484);
  IV  NOT_5179(g3069,I6277);
  IV  NOT_5180(I13776,g8513);
  IV  NOT_5181(I13785,g8516);
  IV  NOT_5182(g1982,g736);
  IV  NOT_5183(g4524,g3946);
  IV  NOT_5184(g6294,I10141);
  IV  NOT_5185(I15500,g10051);
  IV  NOT_5186(I5251,g1424);
  IV  NOT_5187(I6590,g3186);
  IV  NOT_5188(g3540,g3307);
  IV  NOT_5189(I7729,g3757);
  IV  NOT_5190(g5887,I9510);
  IV  NOT_5191(g10356,I15832);
  IV  NOT_5192(I5047,g1185);
  IV  NOT_5193(g5122,g4682);
  IV  NOT_5194(g11500,I17519);
  IV  NOT_5195(g6190,g5426);
  IV  NOT_5196(g2074,g1377);
  IV  NOT_5197(g4319,g4144);
  IV  NOT_5198(g7693,I12326);
  IV  NOT_5199(g11049,I16808);
  IV  NOT_5200(I11950,g6906);
  IV  NOT_5201(I16514,g10717);
  IV  NOT_5202(g10826,I16540);
  IV  NOT_5203(I9062,g4759);
  IV  NOT_5204(g7334,I11650);
  IV  NOT_5205(g10380,I15864);
  IV  NOT_5206(g3206,g2055);
  IV  NOT_5207(I13825,g8488);
  IV  NOT_5208(I13370,g8128);
  IV  NOT_5209(I9620,g5189);
  IV  NOT_5210(g4258,I7509);
  IV  NOT_5211(I16507,g10712);
  IV  NOT_5212(g4352,I7633);
  IV  NOT_5213(I11858,g6888);
  IV  NOT_5214(g11048,I16805);
  IV  NOT_5215(g4577,I7984);
  IV  NOT_5216(g4867,I8204);
  IV  NOT_5217(I14709,g9267);
  IV  NOT_5218(g5033,I8406);
  IV  NOT_5219(g10233,g10187);
  IV  NOT_5220(g6156,g5426);
  IV  NOT_5221(g4717,g3829);
  IV  NOT_5222(I7014,g2919);
  IV  NOT_5223(I12511,g7733);
  IV  NOT_5224(g10182,I15530);
  IV  NOT_5225(g7555,I11989);
  IV  NOT_5226(g7804,I12577);
  IV  NOT_5227(I7414,g4156);
  IV  NOT_5228(I10087,g5753);
  IV  NOT_5229(g9919,I15114);
  IV  NOT_5230(g2080,I4894);
  IV  NOT_5231(I7946,g3417);
  IV  NOT_5232(I10258,g6134);
  IV  NOT_5233(I14087,g8770);
  IV  NOT_5234(g7792,I12541);
  IV  NOT_5235(g2480,I5561);
  IV  NOT_5236(I11367,g6392);
  IV  NOT_5237(I11394,g6621);
  IV  NOT_5238(g5096,g4840);
  IV  NOT_5239(g6942,I11076);
  IV  NOT_5240(g8890,I14236);
  IV  NOT_5241(g2713,g2042);
  IV  NOT_5242(I13367,g8221);
  IV  NOT_5243(I13394,g8137);
  IV  NOT_5244(g4211,I7450);
  IV  NOT_5245(g4186,I7375);
  IV  NOT_5246(g6704,g5949);
  IV  NOT_5247(I17687,g11610);
  IV  NOT_5248(g4386,I7713);
  IV  NOT_5249(g10932,g10827);
  IV  NOT_5250(I8929,g4582);
  IV  NOT_5251(g5845,g5320);
  IV  NOT_5252(g4975,I8351);
  IV  NOT_5253(g2569,I5695);
  IV  NOT_5254(I7513,g4144);
  IV  NOT_5255(g8011,I12853);
  IV  NOT_5256(I17752,g11645);
  IV  NOT_5257(g5195,g4453);
  IV  NOT_5258(g5395,I8831);
  IV  NOT_5259(g5891,g5361);
  IV  NOT_5260(I9842,g5405);
  IV  NOT_5261(I17374,g11411);
  IV  NOT_5262(g7113,I11348);
  IV  NOT_5263(g11106,g10974);
  IV  NOT_5264(g7313,I11587);
  IV  NOT_5265(I11420,g6417);
  IV  NOT_5266(g4426,g3914);
  IV  NOT_5267(g10897,g10827);
  IV  NOT_5268(I12916,g7849);
  IV  NOT_5269(I10069,g5787);
  IV  NOT_5270(g6954,I11100);
  IV  NOT_5271(g6250,I10009);
  IV  NOT_5272(g4170,g3328);
  IV  NOT_5273(g6810,I10840);
  IV  NOT_5274(g4614,g3829);
  IV  NOT_5275(g9527,I14668);
  IV  NOT_5276(g4370,I7671);
  IV  NOT_5277(I12550,g7675);
  IV  NOT_5278(I7378,g4067);
  IV  NOT_5279(I10810,g6539);
  IV  NOT_5280(I11318,g6488);
  IV  NOT_5281(g4125,I7272);
  IV  NOT_5282(I15371,g9990);
  IV  NOT_5283(g6432,g6146);
  IV  NOT_5284(g7908,g7454);
  IV  NOT_5285(I13227,g8264);
  IV  NOT_5286(g6053,I9684);
  IV  NOT_5287(I14955,g9765);
  IV  NOT_5288(I17669,g11604);
  IV  NOT_5289(g8992,I14397);
  IV  NOT_5290(g9764,g9432);
  IV  NOT_5291(I16920,g11084);
  IV  NOT_5292(g11033,I16760);
  IV  NOT_5293(g3291,g2161);
  IV  NOT_5294(I12307,g7245);
  IV  NOT_5295(I5935,g2174);
  IV  NOT_5296(I6844,g2915);
  IV  NOT_5297(g6453,g5817);
  IV  NOT_5298(I9854,g5557);
  IV  NOT_5299(I14970,g9732);
  IV  NOT_5300(g4280,g4013);
  IV  NOT_5301(I7182,g2645);
  IV  NOT_5302(I7288,g2873);
  IV  NOT_5303(g4939,I8303);
  IV  NOT_5304(I11540,g6877);
  IV  NOT_5305(I5982,g2510);
  IV  NOT_5306(g3144,g2462);
  IV  NOT_5307(I11058,g6641);
  IV  NOT_5308(I15795,g10280);
  IV  NOT_5309(g3344,I6528);
  IV  NOT_5310(I16121,g10396);
  IV  NOT_5311(g6568,g5797);
  IV  NOT_5312(I10171,g5992);
  IV  NOT_5313(g4083,I7216);
  IV  NOT_5314(g8080,I12942);
  IV  NOT_5315(I4879,g256);
  IV  NOT_5316(g4544,g3880);
  IV  NOT_5317(g3207,g2439);
  IV  NOT_5318(g8573,I13812);
  IV  NOT_5319(I7916,g3664);
  IV  NOT_5320(I7022,g2941);
  IV  NOT_5321(I13203,g8196);
  IV  NOT_5322(g8480,I13682);
  IV  NOT_5323(g7776,I12493);
  IV  NOT_5324(g2000,g810);
  IV  NOT_5325(I7749,g3764);
  IV  NOT_5326(I6557,g3086);
  IV  NOT_5327(g8713,g8684);
  IV  NOT_5328(I17525,g11486);
  IV  NOT_5329(g2126,g12);
  IV  NOT_5330(g4636,I8036);
  IV  NOT_5331(I15514,g10122);
  IV  NOT_5332(I17424,g11424);
  IV  NOT_5333(g3694,I6851);
  IV  NOT_5334(g6157,I9880);
  IV  NOT_5335(I6071,g2269);
  IV  NOT_5336(I14967,g9763);
  IV  NOT_5337(I12773,g7581);
  IV  NOT_5338(I16682,g10799);
  IV  NOT_5339(I17558,g11504);
  IV  NOT_5340(I15507,g10047);
  IV  NOT_5341(g5081,I8449);
  IV  NOT_5342(I12942,g7982);
  IV  NOT_5343(g3088,I6294);
  IV  NOT_5344(g5815,I9421);
  IV  NOT_5345(g8569,I13800);
  IV  NOT_5346(g4306,g3586);
  IV  NOT_5347(g7965,I12759);
  IV  NOT_5348(I12268,g7107);
  IV  NOT_5349(g5481,I8900);
  IV  NOT_5350(g11507,I17540);
  IV  NOT_5351(I12156,g6878);
  IV  NOT_5352(g4790,g3337);
  IV  NOT_5353(I12655,g7402);
  IV  NOT_5354(g5692,I9221);
  IV  NOT_5355(I15421,g10083);
  IV  NOT_5356(g1964,g114);
  IV  NOT_5357(g10387,g10357);
  IV  NOT_5358(g97,I4780);
  IV  NOT_5359(g7264,I11501);
  IV  NOT_5360(I12180,g7263);
  IV  NOT_5361(g10620,I16295);
  IV  NOT_5362(g4187,I7378);
  IV  NOT_5363(g4061,I7182);
  IV  NOT_5364(g10148,g10121);
  IV  NOT_5365(g11421,I17318);
  IV  NOT_5366(g4387,I7716);
  IV  NOT_5367(g4461,g3829);
  IV  NOT_5368(I6955,g2871);
  IV  NOT_5369(g7360,I11728);
  IV  NOT_5370(g11163,I16920);
  IV  NOT_5371(g10104,I15338);
  IV  NOT_5372(I11146,g6439);
  IV  NOT_5373(g4756,g3440);
  IV  NOT_5374(I17713,g11621);
  IV  NOT_5375(I13738,g8295);
  IV  NOT_5376(I13645,g8379);
  IV  NOT_5377(g8688,g8507);
  IV  NOT_5378(I12335,g7133);
  IV  NOT_5379(g7521,I11901);
  IV  NOT_5380(g10343,I15795);
  IV  NOT_5381(I14010,g8642);
  IV  NOT_5382(I14918,g9535);
  IV  NOT_5383(g8976,I14349);
  IV  NOT_5384(g2608,I5725);
  IV  NOT_5385(I9829,g5013);
  IV  NOT_5386(I16760,g10888);
  IV  NOT_5387(g2220,g104);
  IV  NOT_5388(g4427,g3638);
  IV  NOT_5389(I12930,g7896);
  IV  NOT_5390(g7450,g7148);
  IV  NOT_5391(I12993,g8044);
  IV  NOT_5392(I15473,g10087);
  IV  NOT_5393(I13290,g8254);
  IV  NOT_5394(g2779,g1974);
  IV  NOT_5395(I6150,g2122);
  IV  NOT_5396(g9987,I15187);
  IV  NOT_5397(g11541,g11519);
  IV  NOT_5398(I17610,g11549);
  IV  NOT_5399(I11698,g7057);
  IV  NOT_5400(g4200,I7417);
  IV  NOT_5401(g9771,g9432);
  IV  NOT_5402(I12694,g7374);
  IV  NOT_5403(I12838,g7682);
  IV  NOT_5404(g11473,I17456);
  IV  NOT_5405(g2023,g1357);
  IV  NOT_5406(I10078,g5729);
  IV  NOT_5407(I17255,g11344);
  IV  NOT_5408(g4514,g3946);
  IV  NOT_5409(I10598,g5874);
  IV  NOT_5410(g5783,I9377);
  IV  NOT_5411(g4003,g3144);
  IV  NOT_5412(g7724,I12357);
  IV  NOT_5413(I15359,g10019);
  IV  NOT_5414(I6409,g2356);
  IV  NOT_5415(g8126,I12989);
  IV  NOT_5416(I7719,g3752);
  IV  NOT_5417(g5112,g4682);
  IV  NOT_5418(g7379,g6863);
  IV  NOT_5419(g5218,I8647);
  IV  NOT_5420(g8326,I13360);
  IV  NOT_5421(I17188,g11313);
  IV  NOT_5422(I17124,g11232);
  IV  NOT_5423(g5267,I8711);
  IV  NOT_5424(I17678,g11607);
  IV  NOT_5425(I11427,g6573);
  IV  NOT_5426(I12487,g7723);
  IV  NOT_5427(I15829,g10203);
  IV  NOT_5428(I13427,g8241);
  IV  NOT_5429(g9892,I15079);
  IV  NOT_5430(I8039,g3506);
  IV  NOT_5431(I7752,g3407);
  IV  NOT_5432(g4763,g3586);
  IV  NOT_5433(I12502,g7726);
  IV  NOT_5434(g4191,I7390);
  IV  NOT_5435(I11632,g6931);
  IV  NOT_5436(g7878,g7479);
  IV  NOT_5437(g10850,I16550);
  IV  NOT_5438(g8760,g8670);
  IV  NOT_5439(g11434,I17353);
  IV  NOT_5440(g4391,g3638);
  IV  NOT_5441(g1989,g770);
  IV  NOT_5442(I10322,g6193);
  IV  NOT_5443(g7289,I11543);
  IV  NOT_5444(g7777,I12496);
  IV  NOT_5445(g7658,I12271);
  IV  NOT_5446(g5401,I8839);
  IV  NOT_5447(g3408,g3108);
  IV  NOT_5448(I10159,g5936);
  IV  NOT_5449(g10133,g10064);
  IV  NOT_5450(g5676,I9185);
  IV  NOT_5451(g2451,g248);
  IV  NOT_5452(I10901,g6620);
  IV  NOT_5453(g4637,I8039);
  IV  NOT_5454(I12279,g7225);
  IV  NOT_5455(I5348,g746);
  IV  NOT_5456(g3336,I6523);
  IV  NOT_5457(I15344,g10025);
  IV  NOT_5458(g6778,g5987);
  IV  NOT_5459(g7882,g7479);
  IV  NOT_5460(g3768,I6979);
  IV  NOT_5461(g10896,I16650);
  IV  NOT_5462(I13403,g8236);
  IV  NOT_5463(g11344,I17155);
  IV  NOT_5464(g4307,g4013);
  IV  NOT_5465(g4536,g3880);
  IV  NOT_5466(g10228,I15604);
  IV  NOT_5467(g4159,I7300);
  IV  NOT_5468(g2346,I5414);
  IV  NOT_5469(g4359,g3880);
  IV  NOT_5470(I12469,g7531);
  IV  NOT_5471(g6735,I10736);
  IV  NOT_5472(g8183,I13102);
  IV  NOT_5473(g8608,g8482);
  IV  NOT_5474(g8924,I14249);
  IV  NOT_5475(g5830,I9446);
  IV  NOT_5476(g7611,I12183);
  IV  NOT_5477(g8220,g7826);
  IV  NOT_5478(I12286,g7231);
  IV  NOT_5479(I14561,g9025);
  IV  NOT_5480(g5727,I9273);
  IV  NOT_5481(g2103,I4961);
  IV  NOT_5482(I8919,g4576);
  IV  NOT_5483(g3943,g2779);
  IV  NOT_5484(I9177,g4904);
  IV  NOT_5485(I7233,g2817);
  IV  NOT_5486(I10144,g5689);
  IV  NOT_5487(g9340,I14525);
  IV  NOT_5488(I14295,g8806);
  IV  NOT_5489(I9377,g5576);
  IV  NOT_5490(I17219,g11292);
  IV  NOT_5491(g7799,I12562);
  IV  NOT_5492(g4757,I8109);
  IV  NOT_5493(I16604,g10786);
  IV  NOT_5494(I7054,g3093);
  IV  NOT_5495(I11572,g6822);
  IV  NOT_5496(g8423,I13583);
  IV  NOT_5497(g6475,g5987);
  IV  NOT_5498(g4416,g3638);
  IV  NOT_5499(g7981,g7624);
  IV  NOT_5500(g6949,I11091);
  IV  NOT_5501(g3228,I6409);
  IV  NOT_5502(g8977,I14352);
  IV  NOT_5503(g2732,I5792);
  IV  NOT_5504(I9287,g5576);
  IV  NOT_5505(g9082,g8892);
  IV  NOT_5506(g10310,I15736);
  IV  NOT_5507(g8588,I13831);
  IV  NOT_5508(g7997,g7697);
  IV  NOT_5509(g2753,I5827);
  IV  NOT_5510(I12601,g7629);
  IV  NOT_5511(g6292,I10135);
  IV  NOT_5512(I11127,g6452);
  IV  NOT_5513(g4315,g3863);
  IV  NOT_5514(g4811,g3661);
  IV  NOT_5515(g2508,g940);
  IV  NOT_5516(g8361,I13463);
  IV  NOT_5517(g10379,I15861);
  IV  NOT_5518(I10966,g6561);
  IV  NOT_5519(g2240,g88);
  IV  NOT_5520(I8004,g3967);
  IV  NOT_5521(g2072,I4876);
  IV  NOT_5522(g3433,I6648);
  IV  NOT_5523(I6921,g2839);
  IV  NOT_5524(I5279,g73);
  IV  NOT_5525(g7332,I11644);
  IV  NOT_5526(g10050,I15269);
  IV  NOT_5527(I9199,g4935);
  IV  NOT_5528(g10378,I15858);
  IV  NOT_5529(I8647,g4219);
  IV  NOT_5530(I9399,g5013);
  IV  NOT_5531(g5624,I9056);
  IV  NOT_5532(g7680,g7148);
  IV  NOT_5533(g11506,I17537);
  IV  NOT_5534(g7353,I11707);
  IV  NOT_5535(g2043,g1801);
  IV  NOT_5536(g6084,I9731);
  IV  NOT_5537(g8327,g8164);
  IV  NOT_5538(I14364,g8952);
  IV  NOT_5539(g4874,I8215);
  IV  NOT_5540(g6039,I9652);
  IV  NOT_5541(g5068,g4840);
  IV  NOT_5542(I11956,g6912);
  IV  NOT_5543(g3096,g2482);
  IV  NOT_5544(I13956,g8451);
  IV  NOT_5545(I13376,g8226);
  IV  NOT_5546(I13385,g8230);
  IV  NOT_5547(I11103,g6667);
  IV  NOT_5548(g3496,I6686);
  IV  NOT_5549(g7744,I12397);
  IV  NOT_5550(I11889,g6898);
  IV  NOT_5551(I17470,g11452);
  IV  NOT_5552(g7802,I12571);
  IV  NOT_5553(I5652,g554);
  IV  NOT_5554(g8146,g8033);
  IV  NOT_5555(I5057,g1961);
  IV  NOT_5556(I11354,g6553);
  IV  NOT_5557(g2116,I5020);
  IV  NOT_5558(g8346,I13418);
  IV  NOT_5559(I5843,g2509);
  IV  NOT_5560(I13354,g8214);
  IV  NOT_5561(I8503,g4445);
  IV  NOT_5562(I5989,g2252);
  IV  NOT_5563(I9510,g5421);
  IV  NOT_5564(I11824,g7246);
  IV  NOT_5565(g2034,g1766);
  IV  NOT_5566(g5677,I9188);
  IV  NOT_5567(g8103,g7994);
  IV  NOT_5568(g3395,I6601);
  IV  NOT_5569(g2434,g1362);
  IV  NOT_5570(g3337,g2745);
  IV  NOT_5571(g3913,g2920);
  IV  NOT_5572(I10289,g6003);
  IV  NOT_5573(I17277,g11390);
  IV  NOT_5574(I12168,g7256);
  IV  NOT_5575(I11671,g7047);
  IV  NOT_5576(g9310,I14503);
  IV  NOT_5577(g6583,I10535);
  IV  NOT_5578(g6702,g5949);
  IV  NOT_5579(g4880,g3638);
  IV  NOT_5580(g5866,g5361);
  IV  NOT_5581(g8696,g8656);
  IV  NOT_5582(I5549,g868);
  IV  NOT_5583(I7029,g2946);
  IV  NOT_5584(I14309,g8813);
  IV  NOT_5585(g2347,g1945);
  IV  NOT_5586(I7429,g3344);
  IV  NOT_5587(g10802,I16510);
  IV  NOT_5588(g5149,I8551);
  IV  NOT_5589(I9144,g5007);
  IV  NOT_5590(I14224,g8794);
  IV  NOT_5591(g6919,g6453);
  IV  NOT_5592(I10308,g6003);
  IV  NOT_5593(I12363,g7187);
  IV  NOT_5594(I7956,g3428);
  IV  NOT_5595(g7901,g7712);
  IV  NOT_5596(g4272,g3586);
  IV  NOT_5597(I8320,g4452);
  IV  NOT_5598(g10730,I16407);
  IV  NOT_5599(I12478,g7560);
  IV  NOT_5600(I12015,g6924);
  IV  NOT_5601(g6276,I10087);
  IV  NOT_5602(g11649,I17749);
  IV  NOT_5603(g9824,I14973);
  IV  NOT_5604(g4243,g3524);
  IV  NOT_5605(g3266,I6436);
  IV  NOT_5606(I9259,g5301);
  IV  NOT_5607(g8240,g7972);
  IV  NOT_5608(g2914,I6091);
  IV  NOT_5609(g5198,I8614);
  IV  NOT_5610(g5747,I9317);
  IV  NOT_5611(I15491,g10093);
  IV  NOT_5612(g2210,g103);
  IV  NOT_5613(g4417,I7757);
  IV  NOT_5614(I10495,g6144);
  IV  NOT_5615(g8472,I13666);
  IV  NOT_5616(g6561,g5773);
  IV  NOT_5617(g11648,I17746);
  IV  NOT_5618(g4935,g4420);
  IV  NOT_5619(g9762,I14903);
  IV  NOT_5620(I17419,g11421);
  IV  NOT_5621(I12556,g7678);
  IV  NOT_5622(I15604,g10148);
  IV  NOT_5623(I10816,g6406);
  IV  NOT_5624(I9923,g5308);
  IV  NOT_5625(g2013,g1101);
  IV  NOT_5626(g8443,I13627);
  IV  NOT_5627(g7600,I12150);
  IV  NOT_5628(I12580,g7540);
  IV  NOT_5629(g7574,g6995);
  IV  NOT_5630(I6085,g2234);
  IV  NOT_5631(g10548,I16209);
  IV  NOT_5632(I17155,g11310);
  IV  NOT_5633(g3142,I6360);
  IV  NOT_5634(g5241,g4386);
  IV  NOT_5635(g6527,I10445);
  IV  NOT_5636(I12223,g7049);
  IV  NOT_5637(g4328,g4130);
  IV  NOT_5638(I14687,g9258);
  IV  NOT_5639(I17170,g11294);
  IV  NOT_5640(I14976,g9670);
  IV  NOT_5641(g8116,I12971);
  IV  NOT_5642(g3255,I6421);
  IV  NOT_5643(I7639,g3722);
  IV  NOT_5644(g8316,I13332);
  IV  NOT_5645(g3815,g3228);
  IV  NOT_5646(I11211,g6527);
  IV  NOT_5647(I10374,g5852);
  IV  NOT_5648(g6764,g5987);
  IV  NOT_5649(I7109,g2970);
  IV  NOT_5650(I5909,g2207);
  IV  NOT_5651(I16534,g10747);
  IV  NOT_5652(I10643,g6026);
  IV  NOT_5653(I11088,g6434);
  IV  NOT_5654(I11024,g6399);
  IV  NOT_5655(g9556,I14701);
  IV  NOT_5656(I16098,g10369);
  IV  NOT_5657(g10317,I15749);
  IV  NOT_5658(g8565,I13788);
  IV  NOT_5659(g2820,I5926);
  IV  NOT_5660(g3097,g2482);
  IV  NOT_5661(I9886,g5286);
  IV  NOT_5662(I6941,g2858);
  IV  NOT_5663(g3726,I6898);
  IV  NOT_5664(g7580,I12056);
  IV  NOT_5665(g6503,I10421);
  IV  NOT_5666(g5644,I9093);
  IV  NOT_5667(I5740,g2341);
  IV  NOT_5668(g6970,I11122);
  IV  NOT_5669(g8347,I13421);
  IV  NOT_5670(I15395,g10058);
  IV  NOT_5671(g2317,g622);
  IV  NOT_5672(I8892,g4554);
  IV  NOT_5673(g10129,I15389);
  IV  NOT_5674(g9930,I15127);
  IV  NOT_5675(I9114,g5603);
  IV  NOT_5676(g6925,I11043);
  IV  NOT_5677(I17194,g11317);
  IV  NOT_5678(I7707,g3370);
  IV  NOT_5679(g11395,I17228);
  IV  NOT_5680(g1962,g27);
  IV  NOT_5681(g10057,I15278);
  IV  NOT_5682(g2601,I5704);
  IV  NOT_5683(g10128,I15386);
  IV  NOT_5684(g5818,g5320);
  IV  NOT_5685(g8697,g8660);
  IV  NOT_5686(I6520,g3186);
  IV  NOT_5687(I14668,g9309);
  IV  NOT_5688(g4213,I7456);
  IV  NOT_5689(g11633,I17713);
  IV  NOT_5690(I11659,g7097);
  IV  NOT_5691(I12186,g7264);
  IV  NOT_5692(g6120,I9813);
  IV  NOT_5693(I10195,g6116);
  IV  NOT_5694(I6031,g2209);
  IV  NOT_5695(I12953,g8024);
  IV  NOT_5696(g10323,I15763);
  IV  NOT_5697(g11191,g11112);
  IV  NOT_5698(g2775,I5862);
  IV  NOT_5699(g7076,I11303);
  IV  NOT_5700(I6812,g3290);
  IV  NOT_5701(g3783,I7009);
  IV  NOT_5702(g7476,g6933);
  IV  NOT_5703(I6958,g2872);
  IV  NOT_5704(g5893,g5106);
  IV  NOT_5705(g6277,I10090);
  IV  NOT_5706(I14525,g9109);
  IV  NOT_5707(I14424,g8945);
  IV  NOT_5708(g3112,g2482);
  IV  NOT_5709(g3267,I6439);
  IV  NOT_5710(g10775,I16461);
  IV  NOT_5711(I16766,g10892);
  IV  NOT_5712(I12936,g7983);
  IV  NOT_5713(I15832,g10206);
  IV  NOT_5714(I8340,g4804);
  IV  NOT_5715(I11296,g6525);
  IV  NOT_5716(g2060,g1380);
  IV  NOT_5717(g6617,g6019);
  IV  NOT_5718(I14558,g9024);
  IV  NOT_5719(g6789,I10789);
  IV  NOT_5720(I17749,g11644);
  IV  NOT_5721(I11644,g6970);
  IV  NOT_5722(I17616,g11561);
  IV  NOT_5723(I16871,g10973);
  IV  NOT_5724(I11338,g6680);
  IV  NOT_5725(I13338,g8210);
  IV  NOT_5726(I9594,g5083);
  IV  NOT_5727(g4166,I7315);
  IV  NOT_5728(g11440,I17371);
  IV  NOT_5729(g4366,I7659);
  IV  NOT_5730(g5426,I8869);
  IV  NOT_5731(I15861,g10339);
  IV  NOT_5732(I16360,g10590);
  IV  NOT_5733(I6911,g2825);
  IV  NOT_5734(I13969,g8451);
  IV  NOT_5735(I7833,g3585);
  IV  NOT_5736(g7285,I11531);
  IV  NOT_5737(g3329,I6504);
  IV  NOT_5738(I15247,g10032);
  IV  NOT_5739(g11573,g11561);
  IV  NOT_5740(I5525,g589);
  IV  NOT_5741(I5710,g2431);
  IV  NOT_5742(g3761,I6962);
  IV  NOT_5743(g5614,I9040);
  IV  NOT_5744(I12762,g7541);
  IV  NOT_5745(I17704,g11618);
  IV  NOT_5746(g4056,I7173);
  IV  NOT_5747(g7500,g6943);
  IV  NOT_5748(I10713,g6003);
  IV  NOT_5749(g8317,I13335);
  IV  NOT_5750(I15389,g10110);
  IV  NOT_5751(g4456,g3375);
  IV  NOT_5752(I14713,g9052);
  IV  NOT_5753(g6299,I10156);
  IV  NOT_5754(g5821,I9433);
  IV  NOT_5755(g3828,g2920);
  IV  NOT_5756(g10697,I16370);
  IV  NOT_5757(g6547,g5893);
  IV  NOT_5758(I13197,g8186);
  IV  NOT_5759(g11389,I17216);
  IV  NOT_5760(g11045,I16796);
  IV  NOT_5761(I6733,g3321);
  IV  NOT_5762(I9065,g4760);
  IV  NOT_5763(I17466,g11447);
  IV  NOT_5764(g8601,g8477);
  IV  NOT_5765(g10261,g10126);
  IV  NOT_5766(g2937,I6106);
  IV  NOT_5767(g3727,I6901);
  IV  NOT_5768(g2079,I4891);
  IV  NOT_5769(g5984,I9602);
  IV  NOT_5770(I10610,g5879);
  IV  NOT_5771(g10880,I16610);
  IV  NOT_5772(I15701,g10236);
  IV  NOT_5773(g4355,I7642);
  IV  NOT_5774(g11388,I17213);
  IV  NOT_5775(g7339,I11665);
  IV  NOT_5776(g2479,g26);
  IV  NOT_5777(I10042,g5723);
  IV  NOT_5778(I15272,g10019);
  IV  NOT_5779(I16629,g10860);
  IV  NOT_5780(g2840,I5960);
  IV  NOT_5781(I10189,g6112);
  IV  NOT_5782(g7024,I11169);
  IV  NOT_5783(I16220,g10502);
  IV  NOT_5784(g2190,I5149);
  IV  NOT_5785(g4260,I7513);
  IV  NOT_5786(g2390,I5475);
  IV  NOT_5787(g7795,I12550);
  IV  NOT_5788(I9433,g5069);
  IV  NOT_5789(I17642,g11579);
  IV  NOT_5790(I10678,g5777);
  IV  NOT_5791(g7737,I12388);
  IV  NOT_5792(g7809,I12592);
  IV  NOT_5793(g3703,g2920);
  IV  NOT_5794(I14188,g8792);
  IV  NOT_5795(I14678,g9265);
  IV  NOT_5796(g5106,I8490);
  IV  NOT_5797(g4463,g3829);
  IV  NOT_5798(I9096,g5568);
  IV  NOT_5799(g2156,I5073);
  IV  NOT_5800(g7672,I12293);
  IV  NOT_5801(I14939,g9454);
  IV  NOT_5802(g2356,I5438);
  IV  NOT_5803(g7077,I11306);
  IV  NOT_5804(g6709,g5949);
  IV  NOT_5805(I17733,g11639);
  IV  NOT_5806(g9814,g9490);
  IV  NOT_5807(g5790,I9388);
  IV  NOT_5808(I9550,g5030);
  IV  NOT_5809(I10030,g5685);
  IV  NOT_5810(g7477,I11869);
  IV  NOT_5811(I10093,g5779);
  IV  NOT_5812(I9845,g5405);
  IV  NOT_5813(g3624,I6767);
  IV  NOT_5814(g6140,I9851);
  IV  NOT_5815(g6340,I10243);
  IV  NOT_5816(I5111,g39);
  IV  NOT_5817(I11581,g6826);
  IV  NOT_5818(I11450,g6488);
  IV  NOT_5819(I12568,g7502);
  IV  NOT_5820(g9350,I14555);
  IV  NOT_5821(g10499,I16124);
  IV  NOT_5822(I5311,g98);
  IV  NOT_5823(g3068,g2303);
  IV  NOT_5824(I13714,g8351);
  IV  NOT_5825(I11315,g6644);
  IV  NOT_5826(g8784,I14087);
  IV  NOT_5827(g2942,I6121);
  IV  NOT_5828(g8739,g8640);
  IV  NOT_5829(I12242,g7089);
  IV  NOT_5830(g4279,I7536);
  IV  NOT_5831(I11707,g7009);
  IV  NOT_5832(g7205,I11433);
  IV  NOT_5833(g9773,g9474);
  IV  NOT_5834(I7086,g3142);
  IV  NOT_5835(I13819,g8488);
  IV  NOT_5836(g11061,g10974);
  IV  NOT_5837(g10498,I16121);
  IV  NOT_5838(g9009,I14405);
  IV  NOT_5839(g6435,I10355);
  IV  NOT_5840(g4167,I7318);
  IV  NOT_5841(g5027,I8396);
  IV  NOT_5842(g6517,I10434);
  IV  NOT_5843(g6082,I9727);
  IV  NOT_5844(I12123,g6861);
  IV  NOT_5845(g4318,g4130);
  IV  NOT_5846(g4367,I7662);
  IV  NOT_5847(I16859,g10911);
  IV  NOT_5848(g4872,I8211);
  IV  NOT_5849(g7634,I12242);
  IV  NOT_5850(I5174,g52);
  IV  NOT_5851(I16950,g11081);
  IV  NOT_5852(g8079,I12939);
  IV  NOT_5853(I16370,g10592);
  IV  NOT_5854(g6482,I10412);
  IV  NOT_5855(I11055,g6419);
  IV  NOT_5856(g10056,I15275);
  IV  NOT_5857(I9807,g5419);
  IV  NOT_5858(g8479,g8319);
  IV  NOT_5859(I7185,g2626);
  IV  NOT_5860(I12751,g7626);
  IV  NOT_5861(g9769,I14918);
  IV  NOT_5862(g4057,I7176);
  IV  NOT_5863(g5904,I9539);
  IV  NOT_5864(g7304,I11560);
  IV  NOT_5865(g5200,g4567);
  IV  NOT_5866(g10080,I15308);
  IV  NOT_5867(g8294,I13236);
  IV  NOT_5868(I13978,g8575);
  IV  NOT_5869(g4457,g3829);
  IV  NOT_5870(g2163,I5092);
  IV  NOT_5871(I8877,g4421);
  IV  NOT_5872(g2363,I5441);
  IV  NOT_5873(I7070,g3138);
  IV  NOT_5874(g5446,I8877);
  IV  NOT_5875(I11590,g6829);
  IV  NOT_5876(I16172,g10498);
  IV  NOT_5877(g4193,I7396);
  IV  NOT_5878(g3716,I6876);
  IV  NOT_5879(g11360,I17185);
  IV  NOT_5880(g4393,I7726);
  IV  NOT_5881(I10837,g6717);
  IV  NOT_5882(g2432,I5513);
  IV  NOT_5883(I12293,g7116);
  IV  NOT_5884(g10271,I15665);
  IV  NOT_5885(I12638,g7708);
  IV  NOT_5886(g11447,I17390);
  IV  NOT_5887(I13741,g8296);
  IV  NOT_5888(I15162,g9958);
  IV  NOT_5889(g4549,I7956);
  IV  NOT_5890(I17555,g11503);
  IV  NOT_5891(I6898,g2964);
  IV  NOT_5892(I12265,g7211);
  IV  NOT_5893(g11162,g10950);
  IV  NOT_5894(g7754,I12427);
  IV  NOT_5895(g10461,I15974);
  IV  NOT_5896(g5191,g4640);
  IV  NOT_5897(g8156,I13051);
  IV  NOT_5898(I9248,g4954);
  IV  NOT_5899(g3747,g3015);
  IV  NOT_5900(I11094,g6657);
  IV  NOT_5901(g1973,g466);
  IV  NOT_5902(g5391,I8827);
  IV  NOT_5903(g8356,I13448);
  IV  NOT_5904(g10342,I15792);
  IV  NOT_5905(g3398,g2896);
  IV  NOT_5906(g6214,g5446);
  IV  NOT_5907(g7273,g6365);
  IV  NOT_5908(I5020,g1176);
  IV  NOT_5909(I6510,g3267);
  IV  NOT_5910(g9993,I15193);
  IV  NOT_5911(g10145,I15437);
  IV  NOT_5912(g10031,I15229);
  IV  NOT_5913(g6110,I9783);
  IV  NOT_5914(g5637,I9074);
  IV  NOT_5915(g6310,I10189);
  IV  NOT_5916(g11629,I17701);
  IV  NOT_5917(g9822,I14967);
  IV  NOT_5918(g10199,g10172);
  IV  NOT_5919(g11451,I17410);
  IV  NOT_5920(g11472,I17453);
  IV  NOT_5921(g7044,I11217);
  IV  NOT_5922(g10887,I16623);
  IV  NOT_5923(g2912,I6085);
  IV  NOT_5924(I13735,g8293);
  IV  NOT_5925(g1969,g456);
  IV  NOT_5926(g4121,I7264);
  IV  NOT_5927(g5107,g4459);
  IV  NOT_5928(g8704,g8667);
  IV  NOT_5929(g4321,g3863);
  IV  NOT_5930(g2157,g1703);
  IV  NOT_5931(g11628,I17698);
  IV  NOT_5932(g10198,I15568);
  IV  NOT_5933(I7131,g2640);
  IV  NOT_5934(I7006,g2912);
  IV  NOT_5935(g7983,I12793);
  IV  NOT_5936(I10201,g5998);
  IV  NOT_5937(g5223,g4640);
  IV  NOT_5938(I11695,g7052);
  IV  NOT_5939(g10528,g10464);
  IV  NOT_5940(g10696,g10621);
  IV  NOT_5941(g4232,I7487);
  IV  NOT_5942(I12835,g7660);
  IV  NOT_5943(I13695,g8363);
  IV  NOT_5944(g10330,I15778);
  IV  NOT_5945(g5858,I9475);
  IV  NOT_5946(g10393,g10317);
  IV  NOT_5947(I10075,g5724);
  IV  NOT_5948(I7766,g3770);
  IV  NOT_5949(g8954,I14315);
  IV  NOT_5950(I16540,g10722);
  IV  NOT_5951(g6236,I9981);
  IV  NOT_5952(I6694,g2749);
  IV  NOT_5953(g7543,I11961);
  IV  NOT_5954(I12586,g7561);
  IV  NOT_5955(g11071,g10913);
  IV  NOT_5956(g8363,I13469);
  IV  NOT_5957(I7487,g3371);
  IV  NOT_5958(I8237,g4295);
  IV  NOT_5959(g5416,I8851);
  IV  NOT_5960(I14494,g8887);
  IV  NOT_5961(g3119,I6347);
  IV  NOT_5962(g10132,g10063);
  IV  NOT_5963(I17519,g11484);
  IV  NOT_5964(g10869,I16577);
  IV  NOT_5965(I6088,g2235);
  IV  NOT_5966(I17176,g11286);
  IV  NOT_5967(I17185,g11311);
  IV  NOT_5968(I10623,g6002);
  IV  NOT_5969(I12442,g7672);
  IV  NOT_5970(I17675,g11606);
  IV  NOT_5971(I17092,g11217);
  IV  NOT_5972(I16203,g10454);
  IV  NOT_5973(g4519,I7920);
  IV  NOT_5974(g5251,g4640);
  IV  NOT_5975(g6590,g5949);
  IV  NOT_5976(g6877,I10963);
  IV  NOT_5977(I4777,g18);
  IV  NOT_5978(g10868,I16574);
  IV  NOT_5979(g5811,I9415);
  IV  NOT_5980(g5642,I9087);
  IV  NOT_5981(g3352,I6538);
  IV  NOT_5982(I9783,g5395);
  IV  NOT_5983(g2626,g2000);
  IV  NOT_5984(g7534,I11942);
  IV  NOT_5985(g7729,I12372);
  IV  NOT_5986(g7961,g7664);
  IV  NOT_5987(g5047,g4354);
  IV  NOT_5988(I13457,g8184);
  IV  NOT_5989(I10984,g6757);
  IV  NOT_5990(g9895,I15088);
  IV  NOT_5991(g6657,I10620);
  IV  NOT_5992(g10161,I15479);
  IV  NOT_5993(g4552,g3880);
  IV  NOT_5994(g4606,g3829);
  IV  NOT_5995(I15858,g10336);
  IV  NOT_5996(g8568,I13797);
  IV  NOT_5997(I8089,g3545);
  IV  NOT_5998(I10352,g6216);
  IV  NOT_5999(g6556,g5747);
  IV  NOT_6000(I14352,g8946);
  IV  NOT_6001(g7927,g7500);
  IV  NOT_6002(I10822,g6584);
  IV  NOT_6003(g5874,I9491);
  IV  NOT_6004(I9001,g4762);
  IV  NOT_6005(g10259,g10141);
  IV  NOT_6006(I14418,g8941);
  IV  NOT_6007(g10708,I16387);
  IV  NOT_6008(I16739,g10856);
  IV  NOT_6009(I12430,g7649);
  IV  NOT_6010(g3186,I6373);
  IV  NOT_6011(g5654,I9123);
  IV  NOT_6012(I12493,g7650);
  IV  NOT_6013(g10471,g10378);
  IV  NOT_6014(g7414,I11794);
  IV  NOT_6015(I9293,g5486);
  IV  NOT_6016(g3386,g3144);
  IV  NOT_6017(g10087,I15314);
  IV  NOT_6018(g8357,I13451);
  IV  NOT_6019(I9129,g4892);
  IV  NOT_6020(g7946,g7416);
  IV  NOT_6021(g10258,g10198);
  IV  NOT_6022(g3975,g3121);
  IV  NOT_6023(I7173,g2644);
  IV  NOT_6024(I9329,g5504);
  IV  NOT_6025(I5973,g2247);
  IV  NOT_6026(g4586,g4089);
  IV  NOT_6027(g11394,I17225);
  IV  NOT_6028(g6464,I10398);
  IV  NOT_6029(g7903,g7446);
  IV  NOT_6030(g2683,g2037);
  IV  NOT_6031(I11689,g7044);
  IV  NOT_6032(I6870,g2852);
  IV  NOT_6033(g3274,I6454);
  IV  NOT_6034(g3426,g3121);
  IV  NOT_6035(g5880,g5361);
  IV  NOT_6036(I12035,g6930);
  IV  NOT_6037(I13280,g8250);
  IV  NOT_6038(g2778,g2276);
  IV  NOT_6039(g10244,g10131);
  IV  NOT_6040(I9727,g5250);
  IV  NOT_6041(I7369,g4051);
  IV  NOT_6042(g3370,I6560);
  IV  NOT_6043(I10589,g5763);
  IV  NOT_6044(I13624,g8320);
  IV  NOT_6045(I14194,g8798);
  IV  NOT_6046(g11420,I17315);
  IV  NOT_6047(g6563,g5783);
  IV  NOT_6048(I7920,g3440);
  IV  NOT_6049(g5272,I8724);
  IV  NOT_6050(g11319,I17116);
  IV  NOT_6051(g7036,g6420);
  IV  NOT_6052(g9085,g8892);
  IV  NOT_6053(g10069,I15296);
  IV  NOT_6054(I7459,g3720);
  IV  NOT_6055(I9221,g5236);
  IV  NOT_6056(g4525,g3880);
  IV  NOT_6057(g7436,g7227);
  IV  NOT_6058(g8626,g8498);
  IV  NOT_6059(g6295,I10144);
  IV  NOT_6060(I12517,g7737);
  IV  NOT_6061(I13102,g7928);
  IV  NOT_6062(g6237,I9984);
  IV  NOT_6063(g11446,I17387);
  IV  NOT_6064(g10774,I16458);
  IV  NOT_6065(I17438,g11444);
  IV  NOT_6066(I10477,g6049);
  IV  NOT_6067(I16366,g10591);
  IV  NOT_6068(g5417,I8854);
  IV  NOT_6069(g2075,I4883);
  IV  NOT_6070(I14477,g8943);
  IV  NOT_6071(g10879,I16607);
  IV  NOT_6072(I16632,g10861);
  IV  NOT_6073(g11059,g10974);
  IV  NOT_6074(g6844,I10904);
  IV  NOT_6075(g7335,I11653);
  IV  NOT_6076(g2475,g192);
  IV  NOT_6077(I14119,g8779);
  IV  NOT_6078(g1988,g766);
  IV  NOT_6079(g3544,g3164);
  IV  NOT_6080(g2949,I6150);
  IV  NOT_6081(g7288,I11540);
  IV  NOT_6082(g11540,g11519);
  IV  NOT_6083(g5982,I9598);
  IV  NOT_6084(g10878,I16604);
  IV  NOT_6085(I7793,g3783);
  IV  NOT_6086(I10864,g6634);
  IV  NOT_6087(g3636,I6815);
  IV  NOT_6088(g5629,I9065);
  IV  NOT_6089(I9953,g5484);
  IV  NOT_6090(g6089,g4977);
  IV  NOT_6091(I12193,g7270);
  IV  NOT_6092(g10171,I15507);
  IV  NOT_6093(g6731,g6001);
  IV  NOT_6094(I9068,g4768);
  IV  NOT_6095(g7805,I12580);
  IV  NOT_6096(I5655,g557);
  IV  NOT_6097(g7916,g7651);
  IV  NOT_6098(g11203,g11112);
  IV  NOT_6099(g5542,I8967);
  IV  NOT_6100(g7022,g6389);
  IV  NOT_6101(g3306,I6477);
  IV  NOT_6102(g2998,g2462);
  IV  NOT_6103(g2646,g1992);
  IV  NOT_6104(g4158,g3304);
  IV  NOT_6105(g7422,I11810);
  IV  NOT_6106(g7749,I12412);
  IV  NOT_6107(I6065,g2226);
  IV  NOT_6108(g6557,g5748);
  IV  NOT_6109(I12165,g6882);
  IV  NOT_6110(I12523,g7421);
  IV  NOT_6111(g10792,I16492);
  IV  NOT_6112(g11044,I16793);
  IV  NOT_6113(g3790,g3228);
  IV  NOT_6114(I15281,g10025);
  IV  NOT_6115(g2084,I4900);
  IV  NOT_6116(g2603,I5710);
  IV  NOT_6117(I8967,g4482);
  IV  NOT_6118(g6705,I10682);
  IV  NOT_6119(g2039,g1781);
  IV  NOT_6120(I9677,g5190);
  IV  NOT_6121(g3387,I6587);
  IV  NOT_6122(I10305,g6180);
  IV  NOT_6123(g5800,I9402);
  IV  NOT_6124(I5410,g901);
  IV  NOT_6125(g3461,I6671);
  IV  NOT_6126(I15377,g10104);
  IV  NOT_6127(g6242,I9995);
  IV  NOT_6128(g2850,I5976);
  IV  NOT_6129(g9431,g9085);
  IV  NOT_6130(g7798,I12559);
  IV  NOT_6131(g11301,I17084);
  IV  NOT_6132(g10459,I15968);
  IV  NOT_6133(g9812,g9490);
  IV  NOT_6134(g3756,g3015);
  IV  NOT_6135(g4587,g3829);
  IV  NOT_6136(I12475,g7545);
  IV  NOT_6137(g11377,I17202);
  IV  NOT_6138(I9866,g5274);
  IV  NOT_6139(g6948,I11088);
  IV  NOT_6140(g3622,I6757);
  IV  NOT_6141(g9958,I15157);
  IV  NOT_6142(g7560,I12012);
  IV  NOT_6143(g4275,g3664);
  IV  NOT_6144(g4311,g4130);
  IV  NOT_6145(g10458,I15965);
  IV  NOT_6146(g8782,I14083);
  IV  NOT_6147(g3427,g3144);
  IV  NOT_6148(I15562,g10098);
  IV  NOT_6149(I9349,g5515);
  IV  NOT_6150(g6955,I11103);
  IV  NOT_6151(I10036,g5701);
  IV  NOT_6152(g4615,I8024);
  IV  NOT_6153(g5213,g4640);
  IV  NOT_6154(g11645,I17739);
  IV  NOT_6155(I10177,g6103);
  IV  NOT_6156(I10560,g5887);
  IV  NOT_6157(I11456,g6440);
  IV  NOT_6158(I14101,g8774);
  IV  NOT_6159(I9848,g5557);
  IV  NOT_6160(I15290,g9984);
  IV  NOT_6161(g6254,I10021);
  IV  NOT_6162(g8475,g8314);
  IV  NOT_6163(g4174,I7339);
  IV  NOT_6164(g6814,I10852);
  IV  NOT_6165(g9765,I14910);
  IV  NOT_6166(I17636,g11577);
  IV  NOT_6167(I15698,g10235);
  IV  NOT_6168(g10545,I16200);
  IV  NOT_6169(g2919,I6102);
  IV  NOT_6170(g7037,I11198);
  IV  NOT_6171(g10079,I15305);
  IV  NOT_6172(g10444,g10325);
  IV  NOT_6173(I9699,g5426);
  IV  NOT_6174(g6150,I9869);
  IV  NOT_6175(I14642,g9088);
  IV  NOT_6176(g7437,I11829);
  IV  NOT_6177(I16784,g10895);
  IV  NOT_6178(I5667,g566);
  IV  NOT_6179(I6395,g2334);
  IV  NOT_6180(I6891,g2962);
  IV  NOT_6181(g8292,I13230);
  IV  NOT_6182(g2952,g2455);
  IV  NOT_6183(I16956,g11096);
  IV  NOT_6184(g3345,I6531);
  IV  NOT_6185(I16376,g10596);
  IV  NOT_6186(I13314,g8260);
  IV  NOT_6187(g4284,g3664);
  IV  NOT_6188(g7579,I12053);
  IV  NOT_6189(g8526,I13735);
  IV  NOT_6190(g10598,I16273);
  IV  NOT_6191(g3763,I6968);
  IV  NOT_6192(I10733,g6099);
  IV  NOT_6193(g4545,I7952);
  IV  NOT_6194(I11076,g6649);
  IV  NOT_6195(I11085,g6433);
  IV  NOT_6196(g3391,g2896);
  IV  NOT_6197(g9733,I14876);
  IV  NOT_6198(I15427,g10088);
  IV  NOT_6199(I16095,g10401);
  IV  NOT_6200(g4180,I7357);
  IV  NOT_6201(g5490,I8911);
  IV  NOT_6202(g9270,I14485);
  IV  NOT_6203(g4380,I7701);
  IV  NOT_6204(g11427,I17334);
  IV  NOT_6205(g5166,g4682);
  IV  NOT_6206(I11596,g6831);
  IV  NOT_6207(g4591,g3829);
  IV  NOT_6208(I15632,g10184);
  IV  NOT_6209(g11366,I17191);
  IV  NOT_6210(g3637,I6818);
  IV  NOT_6211(I7216,g2952);
  IV  NOT_6212(g7752,I12421);
  IV  NOT_6213(g11632,I17710);
  IV  NOT_6214(g8484,g8336);
  IV  NOT_6215(I16181,g10491);
  IV  NOT_6216(I10630,g5889);
  IV  NOT_6217(g8439,I13615);
  IV  NOT_6218(g2004,I4820);
  IV  NOT_6219(I10693,g6068);
  IV  NOT_6220(g6836,I10888);
  IV  NOT_6221(I12372,g7137);
  IV  NOT_6222(g7917,g7497);
  IV  NOT_6223(g2986,I6220);
  IV  NOT_6224(g3307,I6480);
  IV  NOT_6225(g9473,g9103);
  IV  NOT_6226(I7671,g3351);
  IV  NOT_6227(g2647,g1993);
  IV  NOT_6228(g10159,I15473);
  IV  NOT_6229(g4420,I7766);
  IV  NOT_6230(g10125,I15377);
  IV  NOT_6231(g10532,g10473);
  IV  NOT_6232(g10901,g10802);
  IV  NOT_6233(I10009,g5542);
  IV  NOT_6234(g5649,I9108);
  IV  NOT_6235(g3359,I6543);
  IV  NOT_6236(I15403,g10069);
  IV  NOT_6237(g1965,g119);
  IV  NOT_6238(g4507,g3546);
  IV  NOT_6239(g5348,I8815);
  IV  NOT_6240(g6967,I11119);
  IV  NOT_6241(I5555,g110);
  IV  NOT_6242(I11269,g6545);
  IV  NOT_6243(g9980,I15181);
  IV  NOT_6244(g2764,I5850);
  IV  NOT_6245(I8462,g4475);
  IV  NOT_6246(g11403,I17252);
  IV  NOT_6247(g10158,I15470);
  IV  NOT_6248(g11547,g11519);
  IV  NOT_6249(g7042,I11211);
  IV  NOT_6250(I11773,g7257);
  IV  NOT_6251(g10783,I16479);
  IV  NOT_6252(g4794,I8164);
  IV  NOT_6253(I11942,g6909);
  IV  NOT_6254(I13773,g8384);
  IV  NOT_6255(I5792,g2080);
  IV  NOT_6256(g7442,g7237);
  IV  NOT_6257(g8702,g8664);
  IV  NOT_6258(I13341,g8210);
  IV  NOT_6259(I12790,g7618);
  IV  NOT_6260(g7786,I12523);
  IV  NOT_6261(g2503,g1872);
  IV  NOT_6262(g3757,I6952);
  IV  NOT_6263(I9352,g4944);
  IV  NOT_6264(I17312,g11392);
  IV  NOT_6265(g10353,I15823);
  IV  NOT_6266(g3416,g3144);
  IV  NOT_6267(g6993,I11135);
  IV  NOT_6268(I11180,g6506);
  IV  NOT_6269(I16190,g10493);
  IV  NOT_6270(I14485,g8883);
  IV  NOT_6271(g7364,I11740);
  IV  NOT_6272(I6815,g2755);
  IV  NOT_6273(I9717,g5426);
  IV  NOT_6274(I15551,g10080);
  IV  NOT_6275(I14555,g9009);
  IV  NOT_6276(g3522,g3164);
  IV  NOT_6277(g8952,I14309);
  IV  NOT_6278(g11572,g11561);
  IV  NOT_6279(I11734,g7024);
  IV  NOT_6280(g8276,I13200);
  IV  NOT_6281(g3811,I7029);
  IV  NOT_6282(g2224,g695);
  IV  NOT_6283(I6097,g2391);
  IV  NOT_6284(g5063,g4363);
  IV  NOT_6285(I10914,g6728);
  IV  NOT_6286(g7454,g7148);
  IV  NOT_6287(I6726,g3306);
  IV  NOT_6288(I14570,g9028);
  IV  NOT_6289(I9893,g5557);
  IV  NOT_6290(I13335,g8206);
  IV  NOT_6291(g7770,I12475);
  IV  NOT_6292(I14914,g9533);
  IV  NOT_6293(g4515,I7916);
  IV  NOT_6294(g4204,I7429);
  IV  NOT_6295(I15127,g9919);
  IV  NOT_6296(I16546,g10724);
  IV  NOT_6297(g8561,I13776);
  IV  NOT_6298(g2320,g18);
  IV  NOT_6299(I10907,g6705);
  IV  NOT_6300(g7725,I12360);
  IV  NOT_6301(I8842,g4556);
  IV  NOT_6302(g7532,I11932);
  IV  NOT_6303(I7308,g3070);
  IV  NOT_6304(g3874,g2920);
  IV  NOT_6305(I8192,g3566);
  IV  NOT_6306(I12208,g7124);
  IV  NOT_6307(I8298,g4437);
  IV  NOT_6308(I8085,g3664);
  IV  NOT_6309(I13965,g8451);
  IV  NOT_6310(g8004,I12838);
  IV  NOT_6311(g6921,I11037);
  IV  NOT_6312(g8986,I14379);
  IV  NOT_6313(I5494,g1690);
  IV  NOT_6314(I13131,g7979);
  IV  NOT_6315(I14239,g8803);
  IV  NOT_6316(I15956,g10402);
  IV  NOT_6317(g2617,g1997);
  IV  NOT_6318(g2906,I6071);
  IV  NOT_6319(I14567,g9027);
  IV  NOT_6320(g2789,g2276);
  IV  NOT_6321(g5619,g4840);
  IV  NOT_6322(g5167,g4682);
  IV  NOT_6323(I15980,g10414);
  AN2 AND2_0(g11103,g2250,g10937);
  AN2 AND2_1(g9900,g9845,g8327);
  AN2 AND2_2(g11095,g845,g10950);
  AN2 AND2_3(g3880,g3186,g2023);
  AN2 AND2_4(g4973,g1645,g4467);
  AN2 AND2_5(g7389,g7001,g3880);
  AN2 AND2_6(g7888,g7465,g7025);
  AN2 AND2_7(g4969,g1642,g4463);
  AN2 AND2_8(g8224,g1882,g7887);
  AN2 AND2_9(g2892,g1980,g1976);
  AN2 AND2_10(g5686,g158,g5361);
  AN2 AND2_11(g10308,g10217,g9085);
  AN2 AND2_12(g4123,g2695,g3037);
  AN2 AND2_13(g8120,g1909,g7944);
  AN2 AND2_14(g6788,g287,g5876);
  AN2 AND2_15(g5598,g778,g4824);
  AN2 AND2_16(g9694,g278,g9432);
  AN2 AND2_17(g10495,g10431,g3971);
  AN2 AND2_18(g2945,g2411,g1684);
  AN2 AND2_19(g11190,g5623,g11065);
  AN2 AND2_20(g8789,g8639,g8719);
  AN2 AND2_21(g9852,g9728,g9563);
  AN2 AND2_22(g5625,g1053,g4399);
  AN2 AND2_23(g4875,g995,g3914);
  AN2 AND2_24(g9701,g1574,g9474);
  AN2 AND2_25(g7138,g6055,g6707);
  AN2 AND2_26(g10752,g10692,g3586);
  AN2 AND2_27(g11211,g11058,g5534);
  AN2 AND2_28(g11024,g435,g10974);
  AN2 AND2_29(g8547,g8307,g7693);
  AN2 AND2_30(g10669,g10577,g9429);
  AN2 AND2_31(g7707,g691,g7206);
  AN2 AND2_32(g4884,g3813,g2971);
  AN2 AND2_33(g4839,g225,g3946);
  AN2 AND2_34(g9870,g1561,g9816);
  AN2 AND2_35(g6640,g5281,g5801);
  AN2 AND2_36(g9650,g2797,g9240);
  AN2 AND2_37(g5687,g139,g5361);
  AN2 AND2_38(g7957,g2885,g7527);
  AN2 AND2_39(g3512,g2050,g2971);
  AN2 AND2_40(g8244,g7847,g4336);
  AN2 AND2_41(g7449,g6868,g4355);
  AN2 AND2_42(g4235,g1011,g3914);
  AN2 AND2_43(g4343,g345,g3586);
  AN2 AND2_44(g11296,g5482,g11241);
  AN2 AND2_45(g9594,g1,g9292);
  AN2 AND2_46(g6829,g213,g6596);
  AN2 AND2_47(g4334,g1160,g3703);
  AN2 AND2_48(g9943,g9923,g9367);
  AN2 AND2_49(g5525,g1721,g4292);
  AN2 AND2_50(g4548,g440,g3990);
  AN3 AND3_0(g8876,g8105,g6764,g8858);
  AN2 AND2_51(g6733,g5678,g4324);
  AN2 AND2_52(g4804,g476,g3458);
  AN2 AND2_53(g10705,g10564,g4840);
  AN2 AND2_54(g9934,g9913,g9624);
  AN2 AND2_55(g6225,g566,g5082);
  AN2 AND2_56(g6324,g1240,g5949);
  AN2 AND2_57(g10686,g10612,g3863);
  AN2 AND2_58(g6540,g1223,g6072);
  AN2 AND2_59(g8663,g8538,g4013);
  AN2 AND2_60(g11581,g1308,g11539);
  AN2 AND2_61(g6206,g560,g5068);
  AN2 AND2_62(g4518,g452,g3975);
  AN2 AND2_63(g3989,g248,g3164);
  AN2 AND2_64(g7730,g7260,g2347);
  AN2 AND2_65(g5174,g1235,g4681);
  AN2 AND2_66(g7504,g7148,g2847);
  AN2 AND2_67(g7185,g1887,g6724);
  AN2 AND2_68(g2563,I5689,I5690);
  AN2 AND2_69(g7881,g7612,g3810);
  AN2 AND2_70(g11070,g2008,g10913);
  AN2 AND2_71(g9859,g9736,g9573);
  AN3 AND3_1(g8877,g8103,g6764,g8858);
  AN2 AND2_72(g11590,g2274,g11561);
  AN2 AND2_73(g6199,g557,g5062);
  AN2 AND2_74(g9266,g8932,g3398);
  AN2 AND2_75(g5545,g1730,g4321);
  AN2 AND2_76(g5180,g4541,g4533);
  AN2 AND2_77(g5591,g1615,g4514);
  AN2 AND2_78(g8556,g8412,g8029);
  AN2 AND2_79(g11094,g374,g10883);
  AN2 AND2_80(g5853,g5044,g1927);
  AN2 AND2_81(g6245,g575,g5098);
  AN2 AND2_82(g4360,g1861,g3748);
  AN3 AND3_2(g8930,g8100,g6368,g8828);
  AN2 AND2_83(g5507,g4310,g3528);
  AN2 AND2_84(g11150,g3087,g10913);
  AN2 AND2_85(g8464,g8302,g7416);
  AN2 AND2_86(g9692,g272,g9432);
  AN2 AND2_87(g4996,g1428,g4682);
  AN2 AND2_88(g7131,g6044,g6700);
  AN2 AND2_89(g11019,g421,g10974);
  AN2 AND2_90(g9960,g9951,g9536);
  AN2 AND2_91(g11196,g4912,g11068);
  AN2 AND2_92(g11018,g7286,g10974);
  AN2 AND2_93(g6819,g243,g6596);
  AN2 AND2_94(g10595,g10550,g4347);
  AN2 AND2_95(g10494,g10433,g3945);
  AN2 AND2_96(g10623,g10544,g4536);
  AN2 AND2_97(g4878,g1868,g3531);
  AN2 AND2_98(g5204,g4838,g2126);
  AN2 AND2_99(g8844,g8609,g8709);
  AN2 AND2_100(g6701,g6185,g4228);
  AN2 AND2_101(g10782,g10725,g5146);
  AN2 AND2_102(g5100,g1791,g4606);
  AN2 AND2_103(g4882,g1089,g3638);
  AN2 AND2_104(g8731,g8622,g7918);
  AN2 AND2_105(g6215,g1504,g5128);
  AN2 AND2_106(g6886,g1932,g6420);
  AN2 AND2_107(g3586,g3323,g2191);
  AN2 AND2_108(g8557,g8415,g8033);
  AN3 AND3_3(g8966,g8081,g6778,g8849);
  AN2 AND2_109(g8071,g691,g7826);
  AN2 AND2_110(g11597,g11576,g5446);
  AN2 AND2_111(g9828,g9722,g9785);
  AN2 AND2_112(g2918,g2411,g1672);
  AN2 AND2_113(g9830,g9725,g9785);
  AN3 AND3_4(g8955,g8110,g6368,g8828);
  AN2 AND2_114(g9592,g4,g9292);
  AN2 AND2_115(g5123,g1618,g4669);
  AN2 AND2_116(g7059,g6078,g6714);
  AN2 AND2_117(g8254,g2773,g7909);
  AN2 AND2_118(g7459,g7148,g2814);
  AN2 AND2_119(g11102,g861,g10950);
  AN2 AND2_120(g7718,g709,g7221);
  AN2 AND2_121(g7535,g7148,g2874);
  AN2 AND2_122(g9703,g1577,g9474);
  AN2 AND2_123(g5528,g4322,g3537);
  AN2 AND2_124(g5151,g4478,g2733);
  AN2 AND2_125(g9932,g9911,g9624);
  AN2 AND2_126(g5530,g1636,g4305);
  AN2 AND2_127(g3506,g986,g2760);
  AN2 AND2_128(g8769,g8629,g5151);
  AN2 AND2_129(g6887,g6187,g6566);
  AN2 AND2_130(g6228,g5605,g713);
  AN2 AND2_131(g6322,g1275,g5949);
  AN2 AND2_132(g3111,I6337,I6338);
  AN3 AND3_5(g8967,g8085,g6778,g8849);
  AN2 AND2_133(g5010,g1458,g4640);
  AN2 AND2_134(g3275,g115,g2356);
  AN2 AND2_135(g10809,g4811,g10754);
  AN2 AND2_136(g2895,g2411,g1678);
  AN2 AND2_137(g7721,g736,g7237);
  AN2 AND2_138(g9866,g1549,g9802);
  AN2 AND2_139(g9716,g1534,g9490);
  AN2 AND2_140(g10808,g10744,g3829);
  AN2 AND2_141(g3374,g1231,g3047);
  AN2 AND2_142(g4492,g1786,g3685);
  AN2 AND2_143(g8822,g8614,g8752);
  AN2 AND2_144(g10560,g10487,g4575);
  AN3 AND3_6(g11456,g3765,g3517,g11422);
  AN2 AND2_145(g9848,g9724,g9557);
  AN2 AND2_146(g4714,g646,g3333);
  AN2 AND2_147(g6550,g1231,g6089);
  AN2 AND2_148(g5172,g4555,g4549);
  AN2 AND2_149(g10642,g10612,g3829);
  AN2 AND2_150(g3284,g2531,g677);
  AN2 AND2_151(g9699,g284,g9432);
  AN2 AND2_152(g9855,g302,g9772);
  AN2 AND2_153(g5618,g1630,g4551);
  AN2 AND2_154(g6891,g1950,g6435);
  AN2 AND2_155(g7940,g7620,g4013);
  AN2 AND2_156(g11085,g312,g10897);
  AN2 AND2_157(g4736,g396,g3379);
  AN2 AND2_158(g4968,g1432,g4682);
  AN2 AND2_159(g8837,g8646,g8697);
  AN2 AND2_160(g9644,g1182,g9125);
  AN2 AND2_161(g5804,g1546,g5261);
  AN2 AND2_162(g8462,g8300,g7406);
  AN4 AND4_0(I6330,g2549,g2556,g2562,g2570);
  AN2 AND2_163(g11156,g333,g10934);
  AN2 AND2_164(g6342,g293,g5886);
  AN2 AND2_165(g9867,g1552,g9807);
  AN2 AND2_166(g9717,g1537,g9490);
  AN2 AND2_167(g4871,g1864,g3523);
  AN2 AND2_168(g10454,g10435,g3411);
  AN2 AND2_169(g4722,g426,g3353);
  AN2 AND2_170(g7741,g6961,g3880);
  AN2 AND2_171(g4500,g1357,g3941);
  AN2 AND2_172(g9386,g1327,g9151);
  AN2 AND2_173(g8842,g8607,g8707);
  AN2 AND2_174(g9599,g8,g9292);
  AN2 AND2_175(g9274,g8974,g5708);
  AN2 AND2_176(g5518,g4317,g3532);
  AN2 AND2_177(g9614,g1197,g9111);
  AN2 AND2_178(g4838,g3275,g4122);
  AN2 AND2_179(g9125,g8966,g6674);
  AN2 AND2_180(g7217,g4610,g6432);
  AN2 AND2_181(g11557,g2707,g11519);
  AN2 AND2_182(g2911,g2411,g1675);
  AN2 AND2_183(g11210,g11078,g4515);
  AN2 AND2_184(g7466,g7148,g2821);
  AN2 AND2_185(g9939,g9918,g9367);
  AN2 AND2_186(g11279,g4939,g11200);
  AN3 AND3_7(g10518,g10513,g10440,I16145);
  AN2 AND2_187(g4477,g1129,g3878);
  AN2 AND2_188(g8708,g7605,g8592);
  AN2 AND2_189(g7055,g5900,g6579);
  AN2 AND2_190(g5264,g1095,g4763);
  AN2 AND2_191(g6329,g1265,g5949);
  AN2 AND2_192(g6828,g1377,g6596);
  AN2 AND2_193(g8176,g5299,g7853);
  AN2 AND2_194(g6830,g1380,g6596);
  AN2 AND2_195(g8005,g7510,g6871);
  AN2 AND2_196(g4099,g770,g3281);
  AN2 AND2_197(g11601,g1351,g11574);
  AN2 AND2_198(g11187,g5597,g11061);
  AN2 AND2_199(g6746,g6228,g6166);
  AN2 AND2_200(g6221,g782,g5598);
  AN2 AND2_201(g8765,g8630,g5151);
  AN2 AND2_202(g9622,g1200,g9111);
  AN2 AND2_203(g11143,g10923,g4567);
  AN2 AND2_204(g9904,g9886,g9676);
  AN2 AND2_205(g8733,g8625,g7920);
  AN3 AND3_8(g8974,g8094,g6368,g8858);
  AN2 AND2_206(g6624,g348,g6171);
  AN2 AND2_207(g11169,g530,g11112);
  AN2 AND2_208(g8073,g709,g7826);
  AN2 AND2_209(g9841,g9706,g9512);
  AN2 AND2_210(g5882,g5592,g3829);
  AN2 AND2_211(g8796,g8645,g8725);
  AN2 AND2_212(g11168,g534,g11112);
  AN2 AND2_213(g4269,g1015,g3914);
  AN2 AND2_214(g5271,g727,g4772);
  AN2 AND2_215(g10348,g10272,g3705);
  AN2 AND2_216(g5611,g1047,g4382);
  AN2 AND2_217(g8069,g673,g7826);
  AN2 AND2_218(g9695,g1567,g9474);
  AN2 AND2_219(g10304,g10211,g9079);
  AN2 AND2_220(g8469,g8305,g7422);
  AN2 AND2_221(g4712,g1071,g3638);
  AN2 AND2_222(g6576,g5762,g5503);
  AN2 AND2_223(g10622,g10543,g4525);
  AN2 AND2_224(g11015,g5217,g10827);
  AN2 AND2_225(g5674,g148,g5361);
  AN2 AND2_226(g9359,g1308,g9173);
  AN2 AND2_227(g9223,g6454,g8960);
  AN2 AND2_228(g11556,g2701,g11519);
  AN2 AND2_229(g9858,g1595,g9774);
  AN2 AND2_230(g5541,g4331,g3582);
  AN2 AND2_231(g4534,g363,g3586);
  AN2 AND2_232(g6198,g1499,g5128);
  AN2 AND2_233(g6747,g2214,g5897);
  AN2 AND2_234(g6699,g6177,g4221);
  AN2 AND2_235(g6855,g1964,g6392);
  AN2 AND2_236(g3804,g3098,g2203);
  AN2 AND2_237(g5680,g153,g5361);
  AN2 AND2_238(g9642,g2654,g9240);
  AN2 AND2_239(g5744,g1528,g5191);
  AN2 AND2_240(g10333,g10262,g3307);
  AN2 AND2_241(g8399,g6094,g8229);
  AN2 AND2_242(g9447,g1762,g9030);
  AN2 AND2_243(g4903,g1849,g4243);
  AN2 AND2_244(g11178,g516,g11112);
  AN2 AND2_245(g8510,g8414,g7972);
  AN2 AND2_246(g8245,g7850,g4339);
  AN2 AND2_247(g6319,g1296,g5949);
  AN2 AND2_248(g11186,g5594,g11059);
  AN2 AND2_249(g3908,g186,g3164);
  AN2 AND2_250(g2951,g2411,g1681);
  AN2 AND2_251(g6352,g278,g5894);
  AN2 AND2_252(g9595,g901,g9205);
  AN2 AND2_253(g4831,g810,g4109);
  AN2 AND2_254(g5492,g1654,g4263);
  AN2 AND2_255(g9272,g8934,g3424);
  AN2 AND2_256(g10312,g10220,g9094);
  AN2 AND2_257(g6186,g546,g5042);
  AN2 AND2_258(g9612,g2652,g9240);
  AN2 AND2_259(g9417,g1738,g9052);
  AN2 AND2_260(g9935,g9914,g9624);
  AN2 AND2_261(g8701,g7597,g8582);
  AN2 AND2_262(g10745,g10658,g3586);
  AN2 AND2_263(g11216,g956,g11162);
  AN2 AND2_264(g9328,g8971,g5708);
  AN2 AND2_265(g11587,g1327,g11546);
  AN2 AND2_266(g6821,g237,g6596);
  AN2 AND2_267(g6325,g1245,g5949);
  AN2 AND2_268(g4560,g431,g4002);
  AN2 AND2_269(g7368,g6980,g3880);
  AN2 AND2_270(g6083,g552,g5619);
  AN2 AND2_271(g6544,g1227,g6081);
  AN2 AND2_272(g5476,g1615,g4237);
  AN2 AND2_273(g7743,g6967,g3880);
  AN2 AND2_274(g4869,g1083,g3638);
  AN2 AND2_275(g5722,g1598,g5144);
  AN2 AND2_276(g6790,g5813,g4398);
  AN2 AND2_277(g8408,g704,g8139);
  AN2 AND2_278(g10761,g10700,g10699);
  AN2 AND2_279(g7734,g6944,g3880);
  AN2 AND2_280(g8136,g7926,g7045);
  AN2 AND2_281(g6187,g5569,g2340);
  AN2 AND2_282(g4752,g401,g3385);
  AN2 AND2_283(g9902,g9894,g9392);
  AN2 AND2_284(g8768,g8623,g5151);
  AN2 AND2_285(g5500,g1657,g4272);
  AN2 AND2_286(g2496,g374,g369);
  AN2 AND2_287(g6756,g3010,g5877);
  AN3 AND3_9(g8972,g8085,g6764,g8858);
  AN2 AND2_288(g6622,g336,g6165);
  AN2 AND2_289(g11639,g11612,g7897);
  AN2 AND2_290(g9366,g1311,g9173);
  AN2 AND2_291(g11230,g471,g11062);
  AN2 AND2_292(g10328,g10252,g3307);
  AN2 AND2_293(g5024,g1284,g4513);
  AN2 AND2_294(g4364,g1215,g3756);
  AN2 AND2_295(g9649,g916,g9205);
  AN2 AND2_296(g5795,g1543,g5251);
  AN2 AND2_297(g5737,g1524,g5183);
  AN2 AND2_298(g6841,g1400,g6596);
  AN2 AND2_299(g4054,g1753,g2793);
  AN2 AND2_300(g6345,g5823,g4426);
  AN2 AND2_301(g11391,g11275,g7912);
  AN2 AND2_302(g9851,g296,g9770);
  AN2 AND2_303(g6763,g5802,g4381);
  AN2 AND2_304(g4770,g416,g3415);
  AN3 AND3_10(I16142,g10511,g10509,g10507);
  AN2 AND2_305(g9698,g1571,g9474);
  AN2 AND2_306(g4725,g1032,g3914);
  AN2 AND2_307(g5477,g1887,g4241);
  AN2 AND2_308(g9964,g9954,g9536);
  AN2 AND2_309(g5523,g1663,g4290);
  AN2 AND2_310(g4553,g435,g3995);
  AN2 AND2_311(g8550,g8402,g8011);
  AN2 AND2_312(g8845,g8611,g8711);
  AN2 AND2_313(g2081,g932,g928);
  AN2 AND2_314(g6359,g281,g5898);
  AN2 AND2_315(g11586,g1324,g11545);
  AN2 AND2_316(g11007,g5147,g10827);
  AN2 AND2_317(g5104,g1796,g4608);
  AN2 AND2_318(g5099,g4821,g3829);
  AN2 AND2_319(g6757,g2221,g5919);
  AN2 AND2_320(g5499,g1627,g4270);
  AN2 AND2_321(g4389,g3529,g3092);
  AN2 AND2_322(g6416,g3497,g5774);
  AN2 AND2_323(g9720,g1546,g9490);
  AN2 AND2_324(g4990,g1444,g4682);
  AN2 AND2_325(g9619,g2772,g9010);
  AN4 AND4_1(I6630,g2677,g2683,g2689,g2701);
  AN2 AND2_326(g6047,g2017,g4977);
  AN2 AND2_327(g9652,g953,g9223);
  AN3 AND3_11(g10515,g10505,g10469,I16142);
  AN2 AND2_328(g9843,g9711,g9519);
  AN2 AND2_329(g5273,g1074,g4776);
  AN2 AND2_330(g11465,g11434,g5446);
  AN2 AND2_331(g5044,g4348,g1918);
  AN2 AND2_332(g11237,g5472,g11109);
  AN2 AND2_333(g9834,g9731,g9785);
  AN2 AND2_334(g6654,g363,g6214);
  AN2 AND2_335(g5444,g1041,g4880);
  AN2 AND2_336(g3714,g1690,g2991);
  AN2 AND2_337(g11340,g11285,g4424);
  AN2 AND2_338(g9598,g2086,g9274);
  AN2 AND2_339(g8097,g6200,g7851);
  AN2 AND2_340(g8726,g8608,g7913);
  AN2 AND2_341(g6880,g4816,g6562);
  AN2 AND2_342(g4338,g1157,g3707);
  AN2 AND2_343(g5543,g4874,g4312);
  AN3 AND3_12(g8960,g8085,g6368,g8828);
  AN2 AND2_344(g4109,g806,g3287);
  AN2 AND2_345(g10759,g10698,g10697);
  AN2 AND2_346(g9938,g9917,g9367);
  AN2 AND2_347(g10758,g10652,g4013);
  AN2 AND2_348(g4759,g406,g3392);
  AN2 AND2_349(g9909,g9891,g9804);
  AN2 AND2_350(g7127,g6663,g2241);
  AN2 AND2_351(g11165,g476,g11112);
  AN2 AND2_352(g6234,g2244,g5151);
  AN2 AND2_353(g6328,g1260,g5949);
  AN2 AND2_354(g8401,g677,g8124);
  AN2 AND2_355(g11006,g5125,g10827);
  AN2 AND2_356(g4865,g1080,g3638);
  AN2 AND2_357(g4715,g1077,g3638);
  AN3 AND3_13(g4604,g3056,g3753,g2325);
  AN2 AND2_358(g5513,g1675,g4282);
  AN2 AND2_359(g11222,g965,g11055);
  AN2 AND2_360(g4498,g1145,g3940);
  AN2 AND2_361(g6554,g5075,g6183);
  AN2 AND2_362(g7732,g6935,g3880);
  AN2 AND2_363(g9586,g2727,g9173);
  AN3 AND3_14(g5178,g2047,g4401,g4104);
  AN2 AND2_364(g4584,g3710,g2322);
  AN2 AND2_365(g7472,g7148,g2829);
  AN2 AND2_366(g11253,g981,g11072);
  AN2 AND2_367(g5182,g1240,g4713);
  AN2 AND2_368(g9860,g1598,g9775);
  AN2 AND2_369(g8703,g7601,g8585);
  AN2 AND2_370(g11600,g1346,g11573);
  AN2 AND2_371(g9710,g1586,g9474);
  AN2 AND2_372(g9645,g1203,g9111);
  AN2 AND2_373(g11236,g5469,g11108);
  AN2 AND2_374(g4162,g3106,g2971);
  AN2 AND2_375(g6090,g553,g5627);
  AN2 AND2_376(g9691,g269,g9432);
  AN2 AND2_377(g11372,g11316,g4266);
  AN2 AND2_378(g6823,g1368,g6596);
  AN2 AND2_379(g11175,g501,g11112);
  AN2 AND2_380(g8068,g664,g7826);
  AN2 AND2_381(g9607,g12,g9274);
  AN2 AND2_382(g9962,g9952,g9536);
  AN2 AND2_383(g6348,g296,g5891);
  AN2 AND2_384(g9659,g956,g9223);
  AN2 AND2_385(g9358,g1318,g9151);
  AN2 AND2_386(g3104,I6316,I6317);
  AN2 AND2_387(g4486,g1711,g3910);
  AN2 AND2_388(g9587,g892,g8995);
  AN2 AND2_389(g5632,g1636,g4563);
  AN2 AND2_390(g9111,g8965,g6674);
  AN2 AND2_391(g4881,g991,g3914);
  AN2 AND2_392(g11209,g11074,g9448);
  AN2 AND2_393(g8848,g8715,g8713);
  AN2 AND2_394(g4070,g3263,g2330);
  AN2 AND2_395(g6463,g5052,g6210);
  AN2 AND2_396(g8699,g7595,g8579);
  AN4 AND4_2(I5689,g1419,g1424,g1428,g1432);
  AN2 AND2_397(g7820,g1896,g7479);
  AN2 AND2_398(g11021,g448,g10974);
  AN2 AND2_399(g5917,g1044,g5320);
  AN2 AND2_400(g6619,g49,g6156);
  AN2 AND2_401(g6318,g1300,g5949);
  AN2 AND2_402(g6872,g1896,g6389);
  AN2 AND2_403(g11320,g11201,g4379);
  AN2 AND2_404(g10514,g10489,g4580);
  AN2 AND2_405(g4006,g201,g3228);
  AN2 AND2_406(g9853,g299,g9771);
  AN2 AND2_407(g11274,g4913,g11197);
  AN2 AND2_408(g6193,g2206,g5151);
  AN2 AND2_409(g8119,g6239,g7890);
  AN2 AND2_410(g9420,g1747,g9030);
  AN2 AND2_411(g5233,g1791,g4492);
  AN2 AND2_412(g7581,g7092,g5420);
  AN2 AND2_413(g6549,g5515,g6175);
  AN2 AND2_414(g11464,g11433,g5446);
  AN2 AND2_415(g4801,g516,g3439);
  AN2 AND2_416(g6834,g1365,g6596);
  AN2 AND2_417(g4487,g1718,g3911);
  AN2 AND2_418(g2939,g2411,g1687);
  AN2 AND2_419(g7060,g6739,g5521);
  AN2 AND2_420(g5770,g4466,g5128);
  AN2 AND2_421(g5725,g1580,g5166);
  AN2 AND2_422(g11641,g11615,g7901);
  AN2 AND2_423(g2544,g1341,g1336);
  AN2 AND2_424(g11292,g11252,g4250);
  AN2 AND2_425(g5532,g1681,g4307);
  AN2 AND2_426(g11153,g3771,g10913);
  AN2 AND2_427(g9905,g9872,g9680);
  AN2 AND2_428(g7739,g6957,g3880);
  AN2 AND2_429(g6321,g1284,g5949);
  AN2 AND2_430(g8386,g6085,g8219);
  AN3 AND3_15(g8975,g8089,g6764,g8858);
  AN2 AND2_431(g2306,g1223,g1218);
  AN2 AND2_432(g6625,g1218,g6178);
  AN2 AND2_433(g7937,g7606,g4013);
  AN2 AND2_434(g10788,g8303,g10754);
  AN2 AND2_435(g10325,g10248,g3307);
  AN2 AND2_436(g8170,g5270,g7853);
  AN2 AND2_437(g5706,g1574,g5121);
  AN2 AND2_438(g2756,g936,g2081);
  AN2 AND2_439(g8821,g8643,g8751);
  AN2 AND2_440(g10946,g5225,g10827);
  AN2 AND2_441(g4169,g2765,g3066);
  AN2 AND2_442(g5029,g1077,g4521);
  AN2 AND2_443(g11164,g4889,g11112);
  AN2 AND2_444(g4007,g2683,g2276);
  AN2 AND2_445(g4059,g1756,g2796);
  AN2 AND2_446(g4868,g1027,g3914);
  AN2 AND2_447(g5675,g131,g5361);
  AN2 AND2_448(g4718,g650,g3343);
  AN2 AND2_449(g10682,g10600,g3863);
  AN2 AND2_450(g6687,g5486,g5840);
  AN2 AND2_451(g7704,g682,g7197);
  AN2 AND2_452(g4582,g525,g4055);
  AN2 AND2_453(g4261,g1019,g3914);
  AN2 AND2_454(g3422,g225,g3228);
  AN2 AND2_455(g5745,g1549,g5192);
  AN2 AND2_456(g8387,g6086,g8220);
  AN2 AND2_457(g7954,g2874,g7512);
  AN2 AND2_458(g11283,g4966,g11205);
  AN2 AND2_459(g8461,g8298,g7403);
  AN2 AND2_460(g10760,g10695,g10691);
  AN2 AND2_461(g11492,g11480,g4807);
  AN3 AND3_16(g7032,g2965,g6626,g5292);
  AN2 AND2_462(g8756,g7431,g8674);
  AN2 AND2_463(g9151,g8967,g6674);
  AN2 AND2_464(g6341,g272,g5885);
  AN2 AND2_465(g10506,g10390,g2135);
  AN2 AND2_466(g9648,g16,g9274);
  AN2 AND2_467(g7453,g7148,g2809);
  AN2 AND2_468(g6525,g5995,g3102);
  AN2 AND2_469(g6645,g67,g6202);
  AN2 AND2_470(g5707,g1595,g5122);
  AN2 AND2_471(g8046,g7548,g5128);
  AN2 AND2_472(g11091,g833,g10950);
  AN2 AND2_473(g11174,g496,g11112);
  AN2 AND2_474(g9010,g6454,g8930);
  AN2 AND2_475(g8403,g6101,g8239);
  AN2 AND2_476(g5201,g1250,g4721);
  AN2 AND2_477(g8841,g8605,g8704);
  AN2 AND2_478(g6879,g1914,g6407);
  AN2 AND2_479(g8763,g7440,g8680);
  AN2 AND2_480(g4502,g2031,g3938);
  AN2 AND2_481(g9839,g9702,g9742);
  AN2 AND2_482(g6358,g5841,g4441);
  AN2 AND2_483(g5575,g1618,g4501);
  AN2 AND2_484(g4940,g3500,g4440);
  AN2 AND2_485(g8107,g6226,g7882);
  AN2 AND2_486(g10240,g10150,g9103);
  AN2 AND2_487(g11192,g5628,g11066);
  AN2 AND2_488(g9618,g910,g9205);
  AN2 AND2_489(g5539,g1684,g4314);
  AN2 AND2_490(g8416,g731,g8151);
  AN2 AND2_491(g9693,g275,g9432);
  AN2 AND2_492(g11553,g2683,g11519);
  AN2 AND2_493(g8047,g7557,g5919);
  AN2 AND2_494(g5268,g1098,g4769);
  AN2 AND2_495(g9555,g9107,g3391);
  AN2 AND2_496(g6180,g2190,g5128);
  AN2 AND2_497(g6832,g1383,g6596);
  AN2 AND2_498(g10633,g10600,g3829);
  AN2 AND2_499(g7894,g7617,g3816);
  AN2 AND2_500(g8654,g8529,g4013);
  AN2 AND2_501(g9621,g1179,g9125);
  AN2 AND2_502(g6794,g5819,g4415);
  AN2 AND2_503(g9313,g8876,g5708);
  AN2 AND2_504(g4883,g248,g3946);
  AN2 AND2_505(g3412,g219,g3228);
  AN2 AND2_506(g7661,g7127,g2251);
  AN3 AND3_17(g2800,g2399,g2369,g591);
  AN2 AND2_507(g3389,g207,g3228);
  AN2 AND2_508(g3706,g471,g3268);
  AN2 AND2_509(g9908,g9890,g9782);
  AN2 AND2_510(g3429,g231,g3228);
  AN2 AND2_511(g6628,g351,g6182);
  AN2 AND2_512(g5470,g1044,g4222);
  AN2 AND2_513(g7526,g7148,g2868);
  AN2 AND2_514(g5897,g2204,g5354);
  AN2 AND2_515(g5025,g1482,g4640);
  AN2 AND2_516(g6204,g3738,g4921);
  AN2 AND2_517(g4048,g1750,g2790);
  AN3 AND3_18(g8935,g8106,g6778,g8849);
  AN2 AND2_518(g3281,g766,g2525);
  AN2 AND2_519(g9593,g898,g9205);
  AN2 AND2_520(g4827,g213,g3946);
  AN2 AND2_521(g10701,g10620,g10619);
  AN2 AND2_522(g10777,g10733,g3015);
  AN2 AND2_523(g8130,g1936,g7952);
  AN2 AND2_524(g9965,g9955,g9536);
  AN2 AND2_525(g3684,g1710,g3015);
  AN2 AND2_526(g11213,g947,g11157);
  AN2 AND2_527(g5006,g1462,g4640);
  AN2 AND2_528(g9933,g9912,g9624);
  AN2 AND2_529(g8554,g8407,g8020);
  AN2 AND2_530(g9641,g913,g9205);
  AN2 AND2_531(g6123,g5630,g4311);
  AN2 AND2_532(g6323,g1235,g5949);
  AN2 AND2_533(g10766,g10646,g4840);
  AN2 AND2_534(g6666,g5301,g5818);
  AN2 AND2_535(g4994,g1504,g4640);
  AN2 AND2_536(g5755,g5103,g5354);
  AN2 AND2_537(g11592,g3717,g11561);
  AN2 AND2_538(g6351,g6210,g5052);
  AN2 AND2_539(g6875,g1905,g6400);
  AN2 AND2_540(g4816,g4070,g2336);
  AN2 AND2_541(g9658,g947,g9240);
  AN2 AND2_542(g6530,g6207,g3829);
  AN2 AND2_543(g8366,g8199,g7265);
  AN2 AND2_544(g9835,g9735,g9785);
  AN2 AND2_545(g6655,g5296,g5812);
  AN3 AND3_19(g5445,g4631,g3875,g2733);
  AN2 AND2_546(g5173,g3094,g4676);
  AN2 AND2_547(g7970,g7384,g7703);
  AN2 AND2_548(g3098,g2331,g2198);
  AN2 AND2_549(g5491,g1624,g4262);
  AN2 AND2_550(g9271,g6681,g8949);
  AN2 AND2_551(g11152,g369,g10903);
  AN2 AND2_552(g9611,g2651,g9010);
  AN2 AND2_553(g6410,g2804,g5759);
  AN2 AND2_554(g10451,g10444,g3365);
  AN2 AND2_555(g4397,g3475,g2181);
  AN2 AND2_556(g7224,g5398,g6441);
  AN2 AND2_557(g5602,g1624,g4535);
  AN2 AND2_558(g4421,g4112,g2980);
  AN2 AND2_559(g6884,g5569,g6564);
  AN2 AND2_560(g6839,g1397,g6596);
  AN2 AND2_561(g8698,g7591,g8576);
  AN3 AND3_20(g8964,g8255,g6368,g8849);
  AN2 AND2_562(g8260,g2775,g7911);
  AN2 AND2_563(g11413,g11354,g10679);
  AN2 AND2_564(g4950,g1415,g4682);
  AN2 AND2_565(g5535,g4327,g3544);
  AN2 AND2_566(g7277,g6772,g731);
  AN2 AND2_567(g8463,g8301,g7410);
  AN2 AND2_568(g3268,g466,g2511);
  AN2 AND2_569(g10785,g10728,g5177);
  AN2 AND2_570(g6618,g658,g6016);
  AN2 AND2_571(g6235,g569,g5089);
  AN2 AND2_572(g10950,g10788,g6355);
  AN2 AND2_573(g4723,g3626,g2779);
  AN2 AND2_574(g8720,g8601,g7905);
  AN2 AND2_575(g6693,g5494,g5845);
  AN2 AND2_576(g11020,g452,g10974);
  AN2 AND2_577(g11583,g1314,g11541);
  AN2 AND2_578(g8118,g1900,g7941);
  AN2 AND2_579(g8167,g5253,g7853);
  AN2 AND2_580(g6334,g1389,g5904);
  AN2 AND2_581(g7892,g7616,g3815);
  AN2 AND2_582(g8652,g8523,g4013);
  AN2 AND2_583(g5721,g1577,g5143);
  AN2 AND2_584(g10367,g10362,g3375);
  AN2 AND2_585(g9901,g9893,g9392);
  AN2 AND2_586(g6792,g290,g5881);
  AN2 AND2_587(g11282,g4958,g11203);
  AN2 AND2_588(g7945,g2847,g7473);
  AN3 AND3_21(g8971,g8081,g6764,g8858);
  AN2 AND2_589(g11302,g5508,g11244);
  AN2 AND2_590(g4585,g521,g4060);
  AN2 AND2_591(g6621,g52,g6164);
  AN2 AND2_592(g5502,g1932,g4275);
  AN2 AND2_593(g11105,g3634,g10937);
  AN2 AND2_594(g7709,g6856,g4333);
  AN2 AND2_595(g8598,g8471,g7432);
  AN2 AND2_596(g7140,g6069,g6711);
  AN2 AND2_597(g9600,g904,g9205);
  AN2 AND2_598(g9864,g1604,g9778);
  AN2 AND2_599(g11640,g11613,g7900);
  AN2 AND2_600(g5188,g4504,g4496);
  AN2 AND2_601(g7435,g7260,g6572);
  AN2 AND2_602(g7876,g7609,g3790);
  AN2 AND2_603(g5030,g1280,g4523);
  AN2 AND2_604(g4058,g2707,g2276);
  AN2 AND2_605(g6776,g5809,g4390);
  AN2 AND2_606(g4890,g630,g4739);
  AN2 AND2_607(g2525,g762,g758);
  AN2 AND2_608(g10301,g8892,g10223);
  AN2 AND2_609(g4505,g354,g3586);
  AN2 AND2_610(g9623,g17,g9274);
  AN2 AND2_611(g10739,g10676,g3368);
  AN2 AND2_612(g11027,g391,g10974);
  AN2 AND2_613(g10738,g10692,g4840);
  AN2 AND2_614(g8687,g8558,g8036);
  AN2 AND2_615(g6360,g302,g5899);
  AN2 AND2_616(g9871,g1564,g9668);
  AN2 AND2_617(g5108,g1801,g4614);
  AN2 AND2_618(g11248,g976,g11071);
  AN2 AND2_619(g4992,g1407,g4682);
  AN2 AND2_620(g11552,g2677,g11519);
  AN2 AND2_621(g9651,g944,g9240);
  AN2 AND2_622(g11204,g971,g11083);
  AN2 AND2_623(g7824,g1932,g7479);
  AN2 AND2_624(g4480,g1133,g3905);
  AN2 AND2_625(g6179,g5115,g5354);
  AN2 AND2_626(g8710,g7607,g8595);
  AN2 AND2_627(g7590,g7102,g5425);
  AN2 AND2_628(g9384,g968,g9223);
  AN2 AND2_629(g3407,g2561,g3012);
  AN2 AND2_630(g9838,g9700,g9754);
  AN2 AND2_631(g3718,g192,g3164);
  AN2 AND2_632(g10661,g10594,g3015);
  AN2 AND2_633(g11380,g11321,g4285);
  AN3 AND3_22(g8879,g8110,g6764,g8858);
  AN2 AND2_634(g7930,g7621,g3110);
  AN3 AND3_23(g8962,g8089,g6368,g8828);
  AN2 AND2_635(g10715,g2272,g10630);
  AN2 AND2_636(g8659,g8535,g4013);
  AN2 AND2_637(g3015,g2028,g2191);
  AN2 AND2_638(g9643,g950,g9223);
  AN2 AND2_639(g9205,g6454,g8957);
  AN2 AND2_640(g5538,g1669,g4313);
  AN2 AND2_641(g4000,g1744,g2778);
  AN2 AND2_642(g4126,g2701,g3040);
  AN2 AND2_643(g4400,g4088,g3829);
  AN2 AND2_644(g2794,I5886,I5887);
  AN2 AND2_645(g4760,g486,g3393);
  AN2 AND2_646(g6238,g572,g5096);
  AN2 AND2_647(g10784,g10727,g5169);
  AN2 AND2_648(g8174,g5284,g7853);
  AN2 AND2_649(g6332,g1374,g5904);
  AN2 AND2_650(g5067,g305,g4811);
  AN2 AND2_651(g5418,g1512,g4344);
  AN2 AND2_652(g10297,g8892,g10211);
  AN2 AND2_653(g6353,g299,g5895);
  AN2 AND2_654(g11026,g386,g10974);
  AN2 AND2_655(g11212,g944,g11155);
  AN2 AND2_656(g6744,g4828,g6151);
  AN2 AND2_657(g5493,g1923,g4265);
  AN2 AND2_658(g10671,g10578,g9431);
  AN2 AND2_659(g4383,g2517,g3829);
  AN2 AND2_660(g5256,g4297,g2779);
  AN2 AND2_661(g4220,g105,g3539);
  AN2 AND2_662(g8380,g8252,g4240);
  AN2 AND2_663(g7071,g5916,g6590);
  AN2 AND2_664(g4779,g501,g3427);
  AN2 AND2_665(g9613,g1176,g9125);
  AN2 AND2_666(g7705,g6853,g4328);
  AN2 AND2_667(g9269,g8933,g3413);
  AN2 AND2_668(g5181,g4520,g4510);
  AN2 AND2_669(g4977,g4567,g4807);
  AN2 AND2_670(g7948,g2855,g7497);
  AN2 AND2_671(g11149,g324,g10930);
  AN2 AND2_672(g9862,g1601,g9777);
  AN2 AND2_673(g11387,g11284,g3629);
  AN2 AND2_674(g7955,g2877,g7516);
  AN2 AND2_675(g4161,g2719,g3060);
  AN2 AND2_676(g11148,g2321,g10913);
  AN2 AND2_677(g9712,g1528,g9490);
  AN2 AND2_678(g8931,g8807,g8164);
  AN2 AND2_679(g11097,g378,g10884);
  AN3 AND3_24(g5421,g4631,g2733,g3819);
  AN2 AND2_680(g11104,g2963,g10937);
  AN2 AND2_681(g5263,g709,g4761);
  AN2 AND2_682(g6092,g1059,g5320);
  AN2 AND2_683(g4999,g1499,g4640);
  AN4 AND4_3(I6338,g2475,g2456,g2451,g2446);
  AN3 AND3_25(g7409,g4976,g632,g6858);
  AN2 AND2_684(g4103,g2683,g2997);
  AN4 AND4_4(I6309,g2446,g2451,g2456,g2475);
  AN2 AND2_685(g6580,g1801,g5944);
  AN2 AND2_686(g5631,g1056,g4416);
  AN2 AND2_687(g9414,g1730,g9052);
  AN2 AND2_688(g9660,g1188,g9125);
  AN2 AND2_689(g9946,g9926,g9392);
  AN2 AND2_690(g5257,g691,g4755);
  AN2 AND2_691(g4732,g391,g3372);
  AN2 AND2_692(g3108,I6330,I6331);
  AN2 AND2_693(g4753,g481,g3386);
  AN2 AND2_694(g9903,g9885,g9673);
  AN2 AND2_695(g10625,g10546,g4552);
  AN2 AND2_696(g5605,g4828,g704);
  AN2 AND2_697(g6623,g55,g6170);
  AN2 AND2_698(g11228,g466,g11060);
  AN2 AND2_699(g11011,g1968,g10809);
  AN2 AND2_700(g6889,g1941,g6427);
  AN2 AND2_701(g8040,g7523,g5128);
  AN2 AND2_702(g7822,g1914,g7479);
  AN2 AND2_703(g8123,g1918,g7946);
  AN2 AND2_704(g11582,g1311,g11540);
  AN2 AND2_705(g4316,g1965,g3400);
  AN2 AND2_706(g10969,g3625,g10809);
  AN2 AND2_707(g5041,g3983,g4401);
  AN2 AND2_708(g9335,g8975,g5708);
  AN2 AND2_709(g9831,g9727,g9785);
  AN2 AND2_710(g4565,g534,g4010);
  AN2 AND2_711(g9422,g1750,g9030);
  AN2 AND2_712(g8648,g4588,g8511);
  AN3 AND3_26(g8875,g8255,g6368,g8858);
  AN2 AND2_713(g5168,g1512,g4679);
  AN2 AND2_714(g7895,g7503,g7036);
  AN2 AND2_715(g8655,g8532,g4013);
  AN2 AND2_716(g3396,g213,g3228);
  AN2 AND2_717(g4914,g1062,g4436);
  AN2 AND2_718(g9947,g9927,g9392);
  AN2 AND2_719(g5772,g1555,g5214);
  AN2 AND2_720(g6838,g192,g6596);
  AN2 AND2_721(g5531,g1666,g4306);
  AN2 AND2_722(g6795,g5036,g5878);
  AN2 AND2_723(g10503,g10388,g2135);
  AN2 AND2_724(g8010,g7738,g7413);
  AN2 AND2_725(g8410,g713,g8143);
  AN2 AND2_726(g6231,g818,g5608);
  AN2 AND2_727(g10581,g10531,g9453);
  AN2 AND2_728(g10450,g10364,g3359);
  AN2 AND2_729(g2804,g2132,g1891);
  AN2 AND2_730(g3418,g2379,g3012);
  AN2 AND2_731(g4820,g186,g3946);
  AN2 AND2_732(g9653,g1185,g9125);
  AN2 AND2_733(g6205,g1515,g5151);
  AN2 AND2_734(g10818,g10730,g4545);
  AN2 AND2_735(g8172,g5275,g7853);
  AN2 AND2_736(g10496,g10429,g3977);
  AN2 AND2_737(g5074,g1771,g4587);
  AN2 AND2_738(g9869,g1558,g9814);
  AN2 AND2_739(g9719,g1543,g9490);
  AN2 AND2_740(g10741,g10635,g4013);
  AN2 AND2_741(g3381,g940,g2756);
  AN2 AND2_742(g5863,g5272,g2173);
  AN2 AND2_743(g8693,g3738,g8509);
  AN2 AND2_744(g5480,g4279,g3519);
  AN2 AND2_745(g4581,g3766,g3254);
  AN2 AND2_746(g3685,g1781,g2981);
  AN2 AND2_747(g5569,g4816,g2338);
  AN2 AND2_748(g8555,g8409,g8025);
  AN2 AND2_749(g3263,g2503,g2328);
  AN2 AND2_750(g9364,g965,g9223);
  AN2 AND2_751(g4784,g506,g3432);
  AN2 AND2_752(g9454,g8994,g5708);
  AN4 AND4_5(I6331,g2060,g2070,g2074,g2077);
  AN2 AND2_753(g11299,g5498,g11243);
  AN2 AND2_754(g6983,g6592,g3105);
  AN2 AND2_755(g7958,g736,g7697);
  AN2 AND2_756(g4995,g1474,g4640);
  AN2 AND2_757(g4079,g2765,g2276);
  AN2 AND2_758(g2264,g1771,g1766);
  AN2 AND2_759(g2160,g745,g746);
  AN2 AND2_760(g3257,g378,g2496);
  AN2 AND2_761(g3101,I6309,I6310);
  AN2 AND2_762(g5000,g1470,g4640);
  AN2 AND2_763(g3301,g1346,g2544);
  AN2 AND2_764(g5126,g3076,g4638);
  AN4 AND4_6(I5084,g1462,g1470,g1474,g1478);
  AN2 AND2_765(g9412,g1727,g9052);
  AN2 AND2_766(g9389,g1330,g9151);
  AN2 AND2_767(g2379,g744,g743);
  AN2 AND2_768(g10706,g10567,g4840);
  AN3 AND3_27(I16145,g10366,g10447,g10446);
  AN2 AND2_769(g10597,g10533,g4359);
  AN3 AND3_28(g8965,g8110,g6778,g8849);
  AN2 AND2_770(g5608,g814,g4831);
  AN2 AND2_771(g5220,g1083,g4729);
  AN2 AND2_772(g10624,g10545,g4544);
  AN2 AND2_773(g10300,g8892,g10220);
  AN2 AND2_774(g5023,g1071,g4511);
  AN2 AND2_775(g4432,g3723,g1975);
  AN2 AND2_776(g4053,g2701,g2276);
  AN2 AND2_777(g8050,g7596,g5919);
  AN2 AND2_778(g5588,g1639,g4508);
  AN3 AND3_29(g6679,g4631,g6074,g2733);
  AN2 AND2_779(g9963,g9953,g9536);
  AN2 AND2_780(g3772,g2542,g3089);
  AN2 AND2_781(g5051,g4432,g2834);
  AN2 AND2_782(g6831,g207,g6596);
  AN2 AND2_783(g2981,g1776,g2264);
  AN2 AND2_784(g8724,g8606,g7910);
  AN2 AND2_785(g4157,g2713,g3055);
  AN2 AND2_786(g9707,g1583,g9474);
  AN3 AND3_30(g8878,g8099,g6368,g8858);
  AN2 AND2_787(g2132,g1872,g1882);
  AN2 AND2_788(g10763,g10639,g4840);
  AN3 AND3_31(g8289,g6777,g8109,g6475);
  AN2 AND2_789(g7898,g7511,g7041);
  AN2 AND2_790(g11271,g5624,g11191);
  AN2 AND2_791(g11461,g11429,g5446);
  AN2 AND2_792(g5732,g1604,g5176);
  AN2 AND2_793(g11145,g315,g10927);
  AN2 AND2_794(g11031,g411,g10974);
  AN2 AND2_795(g9865,g1607,g9780);
  AN2 AND2_796(g5944,g1796,g5233);
  AN2 AND2_797(g9715,g1531,g9490);
  AN2 AND2_798(g9604,g1194,g9111);
  AN2 AND2_799(g8799,g8647,g8727);
  AN2 AND2_800(g11198,g4919,g11069);
  AN2 AND2_801(g6873,g3263,g6557);
  AN2 AND2_802(g6632,g61,g6190);
  AN2 AND2_803(g6095,g1062,g5320);
  AN2 AND2_804(g3863,g3323,g2728);
  AN2 AND2_805(g9833,g9729,g9785);
  AN2 AND2_806(g6653,g70,g6213);
  AN2 AND2_807(g6102,g1038,g5320);
  AN2 AND2_808(g7819,g1887,g7479);
  AN2 AND2_809(g11393,g11280,g7916);
  AN2 AND2_810(g2511,g461,g456);
  AN2 AND2_811(g7088,g2331,g6737);
  AN2 AND2_812(g9584,g2726,g9173);
  AN2 AND2_813(g9896,g9883,g9624);
  AN3 AND3_32(g8209,g4094,g3792,g7980);
  AN2 AND2_814(g6752,g6187,g2343);
  AN2 AND2_815(g4778,g421,g3426);
  AN2 AND2_816(g11161,g1969,g10937);
  AN2 AND2_817(g9268,g6681,g8947);
  AN2 AND2_818(g5681,g135,g5361);
  AN2 AND2_819(g7951,g2868,g7505);
  AN2 AND2_820(g9419,g1744,g9030);
  AN2 AND2_821(g10268,g10183,g3307);
  AN2 AND2_822(g5533,g1724,g4308);
  AN2 AND2_823(g9052,g8936,g7192);
  AN2 AND2_824(g6786,g178,g5919);
  AN2 AND2_825(g10670,g10571,g9091);
  AN2 AND2_826(g11087,g829,g10950);
  AN2 AND2_827(g4949,g3505,g4449);
  AN2 AND2_828(g6364,g5851,g4454);
  AN2 AND2_829(g7825,g1941,g7479);
  AN2 AND2_830(g3400,g115,g3164);
  AN2 AND2_831(g4998,g1304,g4485);
  AN2 AND2_832(g10667,g10576,g9427);
  AN2 AND2_833(g7136,g6050,g6704);
  AN2 AND2_834(g6532,g339,g6057);
  AN2 AND2_835(g9385,g1324,g9151);
  AN4 AND4_7(I5690,g1436,g1440,g1444,g1448);
  AN2 AND2_836(g4484,g1137,g3909);
  AN2 AND2_837(g9897,g9884,g9624);
  AN2 AND2_838(g9425,g1753,g9030);
  AN2 AND2_839(g3383,g186,g3228);
  AN2 AND2_840(g5601,g1035,g4375);
  AN2 AND2_841(g7943,g2840,g7467);
  AN2 AND2_842(g11171,g481,g11112);
  AN2 AND2_843(g3423,I6630,I6631);
  AN2 AND2_844(g7230,g6064,g6444);
  AN2 AND2_845(g4952,g1648,g4457);
  AN2 AND2_846(g8736,g7439,g8635);
  AN2 AND2_847(g6787,g266,g5875);
  AN3 AND3_33(g8968,g8089,g6778,g8849);
  AN2 AND2_848(g10306,g10214,g9082);
  AN2 AND2_849(g9331,g8972,g5708);
  AN2 AND2_850(g11459,g11427,g5446);
  AN2 AND2_851(g4561,g538,g4003);
  AN2 AND2_852(g11425,g11350,g10899);
  AN2 AND2_853(g11458,g11426,g5446);
  AN2 AND2_854(g5739,g1607,g5185);
  AN2 AND2_855(g7496,g7148,g2840);
  AN2 AND2_856(g4986,g1411,g4682);
  AN2 AND2_857(g11010,g5187,g10827);
  AN2 AND2_858(g3999,g1741,g2777);
  AN2 AND2_859(g8175,g5291,g7853);
  AN2 AND2_860(g8722,g8604,g7908);
  AN2 AND2_861(g4764,g411,g3404);
  AN2 AND2_862(g7137,g5590,g6361);
  AN2 AND2_863(g7891,g7471,g7028);
  AN2 AND2_864(g8651,g8520,g4013);
  AN2 AND2_865(g5479,g1845,g4243);
  AN2 AND2_866(g11599,g1341,g11572);
  AN2 AND2_867(g6684,g5314,g5836);
  AN2 AND2_868(g6745,g5605,g6158);
  AN2 AND2_869(g6639,g357,g6196);
  AN2 AND2_870(g10937,g4822,g10822);
  AN2 AND2_871(g3696,g1713,g3015);
  AN2 AND2_872(g4503,g654,g3943);
  AN2 AND2_873(g6791,g269,g5880);
  AN2 AND2_874(g5190,g1245,g4716);
  AN2 AND2_875(g5390,g3220,g4819);
  AN2 AND2_876(g8384,g8180,g3397);
  AN2 AND2_877(g4224,g1092,g3638);
  AN2 AND2_878(g5501,g1672,g4273);
  AN2 AND2_879(g9173,g8968,g6674);
  AN2 AND2_880(g6759,g148,g5919);
  AN2 AND2_881(g8838,g8602,g8702);
  AN2 AND2_882(g8024,g7394,g4337);
  AN2 AND2_883(g10666,g10575,g9424);
  AN2 AND2_884(g11158,g309,g10935);
  AN2 AND2_885(g9602,g2650,g9010);
  AN2 AND2_886(g5704,g143,g5361);
  AN2 AND2_887(g4617,g3275,g3879);
  AN2 AND2_888(g11561,g11518,g3015);
  AN2 AND2_889(g9868,g1555,g9812);
  AN2 AND2_890(g11295,g5475,g11239);
  AN2 AND2_891(g11144,g305,g10926);
  AN2 AND2_892(g9718,g1540,g9490);
  AN2 AND2_893(g3434,g237,g3228);
  AN2 AND2_894(g4987,g1440,g4682);
  AN2 AND2_895(g4771,g496,g3416);
  AN2 AND2_896(g5250,g1270,g4748);
  AN2 AND2_897(g6098,g1065,g5320);
  AN2 AND2_898(g9582,g2725,g9173);
  AN2 AND2_899(g6833,g186,g6596);
  AN2 AND2_900(g3533,g1981,g2892);
  AN2 AND2_901(g4892,g632,g4739);
  AN2 AND2_902(g8104,g6218,g7880);
  AN2 AND2_903(g9415,g1733,g9052);
  AN2 AND2_904(g8499,g8377,g4737);
  AN2 AND2_905(g9664,g1191,g9125);
  AN2 AND2_906(g10740,g10676,g3384);
  AN2 AND2_907(g2534,g798,g794);
  AN2 AND2_908(g8754,g7420,g8667);
  AN2 AND2_909(g9721,g9413,g4785);
  AN2 AND2_910(g6162,g3584,g5200);
  AN2 AND2_911(g4991,g1508,g4640);
  AN2 AND2_912(g6362,g5846,g4450);
  AN4 AND4_8(I6631,g2707,g2713,g2719,g2765);
  AN2 AND2_913(g10685,g10608,g3863);
  AN2 AND2_914(g4340,g1153,g3715);
  AN2 AND2_915(g11023,g440,g10974);
  AN2 AND2_916(g8044,g7598,g5919);
  AN2 AND2_917(g11224,g968,g11056);
  AN2 AND2_918(g11571,g2018,g11561);
  AN2 AND2_919(g4959,g1520,g4682);
  AN2 AND2_920(g10334,g10265,g3307);
  AN2 AND2_921(g5626,g1633,g4557);
  AN2 AND2_922(g9940,g9920,g9367);
  AN2 AND2_923(g4876,g1086,g3638);
  AN2 AND2_924(g6728,g6250,g4318);
  AN2 AND2_925(g6730,g1872,g6128);
  AN2 AND2_926(g9689,g263,g9432);
  AN2 AND2_927(g10762,g10635,g4840);
  AN2 AND2_928(g6070,g1050,g5320);
  AN2 AND2_929(g9428,g1756,g9030);
  AN2 AND2_930(g9030,g8935,g7192);
  AN2 AND2_931(g9430,g1759,g9030);
  AN2 AND2_932(g8927,g7872,g8807);
  AN2 AND2_933(g7068,g5912,g6586);
  AN2 AND2_934(g8014,g7740,g7419);
  AN2 AND2_935(g11392,g11278,g7914);
  AN2 AND2_936(g5782,g1558,g5223);
  AN2 AND2_937(g9910,g9892,g9809);
  AN2 AND2_938(g4824,g774,g4099);
  AN2 AND2_939(g6331,g201,g5904);
  AN2 AND2_940(g4236,g1098,g3638);
  AN2 AND2_941(g11559,g2719,g11519);
  AN2 AND2_942(g9609,g907,g9205);
  AN2 AND2_943(g11558,g2713,g11519);
  AN2 AND2_944(g6087,g1056,g5320);
  AN2 AND2_945(g4877,g243,g3946);
  AN2 AND2_946(g5526,g1950,g4294);
  AN2 AND2_947(g10751,g10646,g4013);
  AN2 AND2_948(g10772,g10655,g4840);
  AN2 AND2_949(g8135,g1945,g7956);
  AN2 AND2_950(g11544,g11515,g10584);
  AN2 AND2_951(g5084,g1776,g4591);
  AN2 AND2_952(g8382,g6077,g8213);
  AN2 AND2_953(g10230,g8892,g10145);
  AN2 AND2_954(g5484,g1896,g4256);
  AN2 AND2_955(g7241,g6772,g6172);
  AN2 AND2_956(g3942,g219,g3164);
  AN2 AND2_957(g10638,g10608,g3829);
  AN2 AND2_958(g4064,g1759,g2799);
  AN2 AND2_959(g9365,g1321,g9151);
  AN2 AND2_960(g9861,g9738,g9579);
  AN2 AND2_961(g8749,g7604,g8660);
  AN2 AND2_962(g11255,g456,g11075);
  AN2 AND2_963(g11189,g5616,g11064);
  AN2 AND2_964(g10510,g10393,g2135);
  AN3 AND3_34(g8947,g8056,g6368,g8828);
  AN2 AND2_965(g2917,g2424,g1657);
  AN2 AND2_966(g5919,g5216,g2965);
  AN2 AND2_967(g11188,g5604,g11063);
  AN2 AND2_968(g9846,g287,g9764);
  AN2 AND2_969(g7818,g1878,g7479);
  AN2 AND2_970(g11460,g11428,g5446);
  AN2 AND2_971(g5276,g736,g4780);
  AN2 AND2_972(g11030,g406,g10974);
  AN2 AND2_973(g11093,g841,g10950);
  AN2 AND2_974(g7893,g7478,g7031);
  AN2 AND2_975(g8653,g8526,g4013);
  AN2 AND2_976(g10442,g10311,g2135);
  AN2 AND2_977(g6535,g345,g6063);
  AN2 AND2_978(g8102,g6209,g7878);
  AN4 AND4_9(I5085,g1490,g1494,g1504,g1508);
  AN2 AND2_979(g5004,g1296,g4499);
  AN2 AND2_980(g3912,g207,g3164);
  AN2 AND2_981(g7186,g2503,g6403);
  AN2 AND2_982(g4489,g348,g3586);
  AN2 AND2_983(g9662,g2094,g9292);
  AN2 AND2_984(g9418,g1741,g9052);
  AN2 AND2_985(g11218,g959,g11053);
  AN2 AND2_986(g4471,g1121,g3862);
  AN2 AND2_987(g10746,g10643,g4013);
  AN2 AND2_988(g7125,g1212,g6648);
  AN2 AND2_989(g7821,g1905,g7479);
  AN2 AND2_990(g6246,g178,g5361);
  AN2 AND2_991(g9256,g6689,g8963);
  AN2 AND2_992(g8042,g7533,g5128);
  AN2 AND2_993(g10237,g10145,g9100);
  AN2 AND2_994(g7939,g2829,g7460);
  AN2 AND2_995(g8786,g8638,g8716);
  AN2 AND2_996(g10684,g10604,g3863);
  AN2 AND2_997(g11455,g11435,g5446);
  AN2 AND2_998(g8364,g658,g8235);
  AN3 AND3_35(g2990,g2061,g2557,g1814);
  AN2 AND2_999(g9847,g290,g9766);
  AN2 AND2_1000(g8054,g7584,g5919);
  AN2 AND2_1001(g5617,g1050,g4391);
  AN2 AND2_1002(g6502,g5981,g3095);
  AN2 AND2_1003(g5789,g1561,g5232);
  AN2 AND2_1004(g4009,g1747,g2789);
  AN2 AND2_1005(g11277,g4920,g11199);
  AN2 AND2_1006(g6940,g6472,g1945);
  AN2 AND2_1007(g7061,g790,g6760);
  AN2 AND2_1008(g11595,g1336,g11575);
  AN2 AND2_1009(g5771,g1534,g5213);
  AN2 AND2_1010(g8553,g8405,g8015);
  AN2 AND2_1011(g4836,g643,g3520);
  AN2 AND2_1012(g5547,g1733,g4326);
  AN2 AND2_1013(g6216,g2232,g5151);
  AN2 AND2_1014(g4967,g1515,g4682);
  AN2 AND2_1015(g6671,g342,g6227);
  AN2 AND2_1016(g7200,g3098,g6418);
  AN2 AND2_1017(g3661,g382,g3257);
  AN2 AND2_1018(g7046,g5892,g6570);
  AN2 AND2_1019(g4229,g999,g3914);
  AN2 AND2_1020(g8389,g6091,g8225);
  AN2 AND2_1021(g6430,g5044,g5791);
  AN2 AND2_1022(g8706,g7602,g8589);
  AN2 AND2_1023(g4993,g1448,g4682);
  AN2 AND2_1024(g6247,g127,g5361);
  AN2 AND2_1025(g9257,g6689,g8964);
  AN2 AND2_1026(g11170,g525,g11112);
  AN2 AND2_1027(g7145,g6082,g6718);
  AN2 AND2_1028(g5738,g1586,g5184);
  AN2 AND2_1029(g6826,g225,g6596);
  AN2 AND2_1030(g7191,g6343,g4323);
  AN2 AND2_1031(g3998,g2677,g2276);
  AN2 AND2_1032(g6741,g3284,g6141);
  AN2 AND2_1033(g5478,g1905,g4242);
  AN2 AND2_1034(g11167,g538,g11112);
  AN2 AND2_1035(g11194,g5637,g11067);
  AN2 AND2_1036(g11589,g1333,g11548);
  AN2 AND2_1037(g6638,g64,g6195);
  AN2 AND2_1038(g4921,g2779,g4431);
  AN2 AND2_1039(g7536,g7148,g2877);
  AN2 AND2_1040(g9585,g889,g8995);
  AN2 AND2_1041(g2957,g2424,g1663);
  AN2 AND2_1042(g11588,g1330,g11547);
  AN2 AND2_1043(g5690,g1567,g5112);
  AN2 AND2_1044(g6883,g1923,g6413);
  AN2 AND2_1045(g4837,g1068,g3638);
  AN3 AND3_36(g8963,g8056,g6368,g8849);
  AN2 AND2_1046(g8791,g8641,g8721);
  AN2 AND2_1047(g6217,g563,g5073);
  AN4 AND4_10(I6316,g2082,g2087,g2381,g2395);
  AN2 AND2_1048(g11022,g444,g10974);
  AN2 AND2_1049(g5915,g4168,g4977);
  AN2 AND2_1050(g4788,g511,g3436);
  AN2 AND2_1051(g8759,g7437,g8677);
  AN2 AND2_1052(g5110,g1806,g4618);
  AN2 AND2_1053(g11254,g986,g11073);
  AN2 AND2_1054(g6827,g219,g6596);
  AN3 AND3_37(g8957,g8081,g6368,g8828);
  AN2 AND2_1055(g6333,g197,g5904);
  AN2 AND2_1056(g8049,g7567,g5919);
  AN2 AND2_1057(g4392,g3273,g3829);
  AN2 AND2_1058(g9856,g1592,g9773);
  AN2 AND2_1059(g9411,g1724,g9052);
  AN2 AND2_1060(g5002,g1494,g4640);
  AN2 AND2_1061(g11101,g857,g10950);
  AN2 AND2_1062(g11177,g511,g11112);
  AN2 AND2_1063(g11560,g2765,g11519);
  AN2 AND2_1064(g8098,g6201,g7852);
  AN2 AND2_1065(g3970,g225,g3164);
  AN2 AND2_1066(g4941,g1038,g4451);
  AN2 AND2_1067(g10453,g10437,g3395);
  AN2 AND2_1068(g5877,g4921,g639);
  AN2 AND2_1069(g6662,g366,g6220);
  AN2 AND2_1070(g7935,g2821,g7454);
  AN2 AND2_1071(g6067,g1047,g5320);
  AN4 AND4_11(I6317,g2406,g2420,g2434,g2438);
  AN2 AND2_1072(g9863,g9740,g9576);
  AN4 AND4_12(I5886,g174,g170,g2249,g2254);
  AN2 AND2_1073(g6994,g6758,g3829);
  AN2 AND2_1074(g9713,g1589,g9474);
  AN2 AND2_1075(g4431,g2268,g3533);
  AN2 AND2_1076(g4252,g1007,g3914);
  AN2 AND2_1077(g11166,g542,g11112);
  AN2 AND2_1078(g7130,g6041,g6697);
  AN2 AND2_1079(g11009,g5179,g10827);
  AN2 AND2_1080(g7542,g7148,g2885);
  AN2 AND2_1081(g8019,g7386,g4332);
  AN2 AND2_1082(g11008,g5171,g10827);
  AN2 AND2_1083(g3516,g1209,g3015);
  AN2 AND2_1084(g8052,g7573,g5128);
  AN2 AND2_1085(g3987,g243,g3164);
  AN2 AND2_1086(g4765,g491,g3405);
  AN2 AND2_1087(g11555,g2695,g11519);
  AN2 AND2_1088(g9857,g9734,g9569);
  AN2 AND2_1089(g8728,g8610,g7915);
  AN2 AND2_1090(g8730,g8613,g7917);
  AN2 AND2_1091(g8185,g664,g7997);
  AN2 AND2_1092(g5194,g1610,g4717);
  AN2 AND2_1093(g8385,g6084,g8218);
  AN2 AND2_1094(g4610,g3804,g2212);
  AN2 AND2_1095(g7902,g7661,g6587);
  AN2 AND2_1096(g4073,g3200,g3222);
  AN2 AND2_1097(g8070,g682,g7826);
  AN2 AND2_1098(g5731,g1583,g5175);
  AN2 AND2_1099(g11238,g5474,g11110);
  AN2 AND2_1100(g4473,g1125,g3874);
  AN2 AND2_1101(g8470,g8308,g7427);
  AN2 AND2_1102(g5489,g4287,g3521);
  AN2 AND2_1103(g3991,g1738,g2774);
  AN4 AND4_13(I5887,g2078,g2083,g166,g2095);
  AN2 AND2_1104(g7823,g1923,g7479);
  AN2 AND2_1105(g4069,g1762,g2802);
  AN3 AND3_38(g11519,g1317,g3015,g11492);
  AN2 AND2_1106(g11176,g506,g11112);
  AN2 AND2_1107(g11092,g837,g10950);
  AN2 AND2_1108(g11154,g330,g10932);
  AN2 AND2_1109(g9608,g7,g9292);
  AN2 AND2_1110(g11637,g11626,g5446);
  AN2 AND2_1111(g2091,g976,g971);
  AN2 AND2_1112(g8406,g695,g8131);
  AN2 AND2_1113(g5254,g4335,g4165);
  AN2 AND2_1114(g7260,g6752,g2345);
  AN2 AND2_1115(g5150,g1275,g4678);
  AN2 AND2_1116(g8766,g8612,g5151);
  AN2 AND2_1117(g9588,g3272,g9173);
  AN2 AND2_1118(g8801,g8742,g8729);
  AN2 AND2_1119(g7063,g5903,g6582);
  AN2 AND2_1120(g10303,g10208,g9076);
  AN2 AND2_1121(g5009,g1486,g4640);
  AN2 AND2_1122(g9665,g1314,g9151);
  AN2 AND2_1123(g8748,g7670,g8656);
  AN2 AND2_1124(g11215,g953,g11160);
  AN2 AND2_1125(g10750,g10687,g3586);
  AN3 AND3_39(g5769,g2112,g4921,g3818);
  AN2 AND2_1126(g8755,g7426,g8671);
  AN2 AND2_1127(g6673,g5305,g5822);
  AN2 AND2_1128(g5212,g1255,g4726);
  AN2 AND2_1129(g7720,g727,g7232);
  AN3 AND3_40(g5918,g2965,g5292,g4609);
  AN2 AND2_1130(g8045,g7547,g5128);
  AN2 AND2_1131(g8173,g7971,g3112);
  AN2 AND2_1132(g11349,g11288,g7964);
  AN2 AND2_1133(g7843,g7599,g5919);
  AN2 AND2_1134(g9696,g281,g9432);
  AN2 AND2_1135(g6772,g6228,g722);
  AN2 AND2_1136(g6058,g1035,g5320);
  AN2 AND2_1137(g6531,g79,g6056);
  AN2 AND2_1138(g6743,g4106,g6146);
  AN2 AND2_1139(g6890,g6752,g6568);
  AN2 AND2_1140(g7549,g7269,g3829);
  AN2 AND2_1141(g8169,g5265,g7853);
  AN2 AND2_1142(g11304,g5520,g11245);
  AN2 AND2_1143(g9944,g9924,g9392);
  AN2 AND2_1144(g9240,g6454,g8962);
  AN2 AND2_1145(g8059,g7592,g5919);
  AN2 AND2_1146(g8718,g8600,g7903);
  AN2 AND2_1147(g8767,g8616,g5151);
  AN2 AND2_1148(g9316,g8877,g5708);
  AN2 AND2_1149(g7625,g673,g7085);
  AN2 AND2_1150(g8793,g8644,g8723);
  AN2 AND2_1151(g2940,g2424,g1654);
  AN2 AND2_1152(g4114,g1351,g3301);
  AN2 AND2_1153(g11636,g11624,g7936);
  AN2 AND2_1154(g10949,g2947,g10809);
  AN2 AND2_1155(g4870,g237,g3946);
  AN2 AND2_1156(g3563,g3275,g2126);
  AN2 AND2_1157(g10948,g2223,g10809);
  AN2 AND2_1158(g8246,g7846,g7442);
  AN2 AND2_1159(g5788,g1540,g5231);
  AN2 AND2_1160(g4008,g2689,g2276);
  AN2 AND2_1161(g9596,g2649,g9010);
  AN2 AND2_1162(g5249,g1089,g4747);
  AN2 AND2_1163(g11585,g1321,g11543);
  AN2 AND2_1164(g3089,g2054,g2050);
  AN2 AND2_1165(g4972,g1436,g4682);
  AN2 AND2_1166(g11554,g2689,g11519);
  AN2 AND2_1167(g7586,g7096,g5423);
  AN2 AND2_1168(g10673,g10580,g9450);
  AN3 AND3_41(g4806,g3215,g3992,g2493);
  AN2 AND2_1169(g5485,g1914,g4257);
  AN2 AND2_1170(g9936,g9915,g9624);
  AN2 AND2_1171(g2910,g2424,g1660);
  AN2 AND2_1172(g9317,g6109,g8875);
  AN2 AND2_1173(g10933,g10853,g3982);
  AN2 AND2_1174(g8388,g8177,g7689);
  AN2 AND2_1175(g4465,g1117,g3828);
  AN2 AND2_1176(g7141,g6073,g6716);
  AN2 AND2_1177(g10508,g10391,g2135);
  AN2 AND2_1178(g4230,g1095,g3638);
  AN2 AND2_1179(g10634,g10604,g3829);
  AN2 AND2_1180(g9601,g922,g9192);
  AN2 AND2_1181(g6126,g5639,g4319);
  AN2 AND2_1182(g6326,g1250,g5949);
  AN2 AND2_1183(g7710,g700,g7214);
  AN2 AND2_1184(g8028,g7375,g7436);
  AN2 AND2_1185(g6760,g786,g6221);
  AN2 AND2_1186(g5640,g1059,g4427);
  AN2 AND2_1187(g5031,g1478,g4640);
  AN2 AND2_1188(g4550,g342,g3586);
  AN2 AND2_1189(g7879,g7610,g3798);
  AN2 AND2_1190(g7962,g7730,g6712);
  AN2 AND2_1191(g9597,g1170,g9125);
  AN2 AND2_1192(g10452,g10439,g3388);
  AN2 AND2_1193(g4891,g631,g4739);
  AN2 AND2_1194(g5005,g1490,g4640);
  AN2 AND2_1195(g6423,g4348,g5784);
  AN2 AND2_1196(g8108,g1891,g7938);
  AN3 AND3_42(g4807,g3015,g1289,g3937);
  AN2 AND2_1197(g5911,g3322,g4977);
  AN2 AND2_1198(g9937,g9916,g9624);
  AN2 AND2_1199(g9840,g9704,g9747);
  AN2 AND2_1200(g10780,g10723,g5124);
  AN2 AND2_1201(g8217,g1872,g7883);
  AN2 AND2_1202(g11013,g5209,g10827);
  AN2 AND2_1203(g9390,g1333,g9151);
  AN2 AND2_1204(g11214,g950,g11159);
  AN2 AND2_1205(g6327,g1255,g5949);
  AN2 AND2_1206(g4342,g1149,g3719);
  AN2 AND2_1207(g5796,g1564,g5252);
  AN2 AND2_1208(g5473,g4268,g3518);
  AN2 AND2_1209(g6346,g5038,g5883);
  AN2 AND2_1210(g6633,g354,g6191);
  AN2 AND2_1211(g11005,g5119,g10827);
  AN2 AND2_1212(g8365,g668,g8240);
  AN2 AND2_1213(g8048,g7558,g5919);
  AN2 AND2_1214(g4481,g1713,g3906);
  AN2 AND2_1215(g4097,g2677,g2989);
  AN2 AND2_1216(g8055,g7588,g5128);
  AN2 AND2_1217(g4497,g351,g3586);
  AN2 AND2_1218(g9942,g9922,g9367);
  AN2 AND2_1219(g6696,g5504,g5850);
  AN3 AND3_43(g10731,g5118,g1850,g10665);
  AN2 AND2_1220(g8827,g8552,g8696);
  AN2 AND2_1221(g5540,g1727,g4315);
  AN2 AND2_1222(g4960,g1403,g4682);
  AN2 AND2_1223(g8846,g8615,g8712);
  AN2 AND2_1224(g6508,g5983,g3096);
  AN2 AND2_1225(g6240,g182,g5361);
  AN2 AND2_1226(g7931,g2809,g7446);
  AN2 AND2_1227(g5287,g3876,g4782);
  AN2 AND2_1228(g6472,g5853,g1936);
  AN2 AND2_1229(g11100,g853,g10950);
  AN2 AND2_1230(g11235,g5443,g11107);
  AN2 AND2_1231(g5199,g1068,g4719);
  AN2 AND2_1232(g6316,g1270,g5949);
  AN2 AND2_1233(g7515,g7148,g2855);
  AN2 AND2_1234(g10583,g10518,g10515);
  AN2 AND2_1235(g5781,g1537,g5222);
  AN2 AND2_1236(g8018,g7742,g7425);
  AN2 AND2_1237(g4401,g2971,g3772);
  AN3 AND3_44(g8994,g8110,g6778,g8925);
  AN2 AND2_1238(g2950,g2424,g1666);
  AN2 AND2_1239(g5510,g1630,g4280);
  AN2 AND2_1240(g6347,g275,g5890);
  AN2 AND2_1241(g9357,g962,g9223);
  AN2 AND2_1242(g4828,g4106,g695);
  AN2 AND2_1243(g11407,g11339,g5949);
  AN2 AND2_1244(g4727,g386,g3364);
  AN2 AND2_1245(g10357,g10278,g2462);
  AN2 AND2_1246(g10743,g10639,g4013);
  AN2 AND2_1247(g5259,g627,g4739);
  AN2 AND2_1248(g5694,g162,g5361);
  AN2 AND2_1249(g10769,g10652,g4840);
  AN2 AND2_1250(g11584,g1318,g11542);
  AN2 AND2_1251(g4932,g1065,g4442);
  AN2 AND2_1252(g10768,g10649,g4840);
  AN2 AND2_1253(g6820,g1362,g6596);
  AN2 AND2_1254(g4068,g2719,g2276);
  AN2 AND2_1255(g6317,g1304,g5949);
  AN2 AND2_1256(g5215,g4276,g3400);
  AN2 AND2_1257(g4576,g530,g4049);
  AN2 AND2_1258(g4866,g231,g3946);
  AN2 AND2_1259(g6775,g822,g6231);
  AN2 AND2_1260(g3829,g2028,g2728);
  AN2 AND2_1261(g10662,g8892,g10571);
  AN2 AND2_1262(g8101,g6208,g7877);
  AN2 AND2_1263(g5825,g3204,g5318);
  AN4 AND4_14(I6310,g2396,g2407,g2421,g2435);
  AN2 AND2_1264(g7884,g7457,g7022);
  AN2 AND2_1265(g5008,g1292,g4507);
  AN2 AND2_1266(g3974,g231,g3164);
  AN2 AND2_1267(g9949,g9929,g9392);
  AN2 AND2_1268(g2531,g658,g668);
  AN2 AND2_1269(g9292,g8878,g5708);
  AN2 AND2_1270(g10778,g1027,g10729);
  AN2 AND2_1271(g8041,g7524,g5128);
  AN2 AND2_1272(g6079,g1053,g5320);
  AN2 AND2_1273(g7235,g6663,g6447);
  AN2 AND2_1274(g9603,g1173,g9125);
  AN2 AND2_1275(g6840,g248,g6596);
  AN2 AND2_1276(g9850,g9726,g9560);
  AN2 AND2_1277(g7988,g1878,g7379);
  AN2 AND2_1278(g5228,g1086,g4734);
  AN2 AND2_1279(g7134,g5587,g6354);
  AN2 AND2_1280(g5934,g5215,g1965);
  AN2 AND2_1281(g5230,g1265,g4735);
  AN2 AND2_1282(g8168,g5262,g7853);
  AN2 AND2_1283(g9583,g886,g8995);
  AN2 AND2_1284(g10672,g10579,g9449);
  AN2 AND2_1285(g3287,g802,g2534);
  AN2 AND2_1286(g8772,g8627,g5151);
  AN2 AND2_1287(g4893,g635,g4739);
  AN2 AND2_1288(g10331,g10256,g3307);
  AN2 AND2_1289(g8505,g8309,g4789);
  AN2 AND2_1290(g10449,g10420,g3345);
  AN2 AND2_1291(g11273,g5638,g11195);
  AN2 AND2_1292(g8734,g8626,g7923);
  AN2 AND2_1293(g5913,g1041,g5320);
  AN2 AND2_1294(g10448,g10421,g3335);
  AN2 AND2_1295(g6163,g4572,g5354);
  AN2 AND2_1296(g6363,g284,g5901);
  AN2 AND2_1297(g7202,g6349,g4329);
  AN2 AND2_1298(g11463,g11432,g5446);
  AN2 AND2_1299(g8074,g718,g7826);
  AN2 AND2_1300(g4325,g1166,g3682);
  AN2 AND2_1301(g8474,g8383,g5285);
  AN2 AND2_1302(g11234,g5424,g11106);
  AN2 AND2_1303(g5266,g718,g4766);
  AN2 AND2_1304(g4483,g336,g3586);
  AN2 AND2_1305(g5248,g673,g4738);
  AN2 AND2_1306(g11514,g11491,g5151);
  AN2 AND2_1307(g5255,g682,g4754);
  AN2 AND2_1308(g4106,g3284,g686);
  AN2 AND2_1309(g2760,g981,g2091);
  AN2 AND2_1310(g5097,g1786,g4603);
  AN2 AND2_1311(g5726,g1601,g5167);
  AN2 AND2_1312(g5497,g4296,g3522);
  AN2 AND2_1313(g5354,g2733,g4460);
  AN2 AND2_1314(g7933,g2814,g7450);
  AN2 AND2_1315(g9617,g9,g9274);
  AN2 AND2_1316(g9906,g9873,g9683);
  AN2 AND2_1317(g11012,g5196,g10827);
  AN2 AND2_1318(g7050,g5896,g6575);
  AN2 AND2_1319(g10971,g10849,g3161);
  AN2 AND2_1320(g4904,g1850,g4243);
  AN2 AND2_1321(g10369,g10361,g3382);
  AN2 AND2_1322(g8400,g6097,g8234);
  AN2 AND2_1323(g4345,g1169,g3730);
  AN2 AND2_1324(g2161,I5084,I5085);
  AN2 AND2_1325(g5001,g1300,g4491);
  AN2 AND2_1326(g9945,g9925,g9392);
  AN2 AND2_1327(g7271,g5028,g6499);
  AN2 AND2_1328(g9709,g1524,g9490);
  AN2 AND2_1329(g4223,g1003,g3914);
  AN2 AND2_1330(g10716,g10497,g10675);
  AN2 AND2_1331(g11291,g11247,g4233);
  AN2 AND2_1332(g6661,g73,g6219);
  AN2 AND2_1333(g11173,g491,g11112);
  AN2 AND2_1334(g6075,g549,g5613);
  AN2 AND2_1335(g8023,g7367,g7430);
  AN2 AND2_1336(g9907,g9888,g9686);
  AN2 AND2_1337(g10582,g10532,g9473);
  AN2 AND2_1338(g5746,g1589,g5193);
  AN2 AND2_1339(g5221,g1260,g4730);
  AN2 AND2_1340(g9959,g9950,g9536);
  AN2 AND2_1341(g7674,g7004,g3880);
  AN2 AND2_1342(g9690,g266,g9432);
  AN2 AND2_1343(g6627,g58,g6181);
  AN2 AND2_1344(g5703,g174,g5361);
  AN2 AND2_1345(g4522,g360,g3586);
  AN2 AND2_1346(g4115,g2689,g3009);
  AN2 AND2_1347(g7541,g7075,g3109);
  AN2 AND2_1348(g10627,g10548,g4564);
  AN2 AND2_1349(g4047,g2695,g2276);
  AN2 AND2_1350(g6526,g76,g6052);
  AN2 AND2_1351(g2944,g2424,g1669);
  AN2 AND2_1352(g6646,g360,g6203);
  AN2 AND2_1353(g7132,g6048,g6702);
  AN2 AND2_1354(g11029,g401,g10974);
  AN2 AND2_1355(g8051,g7572,g5128);
  AN2 AND2_1356(g8127,g1927,g7949);
  AN2 AND2_1357(g7209,g3804,g6425);
  AN2 AND2_1358(g11028,g396,g10974);
  AN2 AND2_1359(g6439,g4479,g5919);
  AN2 AND2_1360(g10742,g10655,g3586);
  AN2 AND2_1361(g9110,g8880,g4790);
  AN2 AND2_1362(g10681,g10567,g3586);
  AN2 AND2_1363(g4537,g444,g3988);
  AN2 AND2_1364(g9663,g959,g9223);
  AN2 AND2_1365(g5349,g2126,g4617);
  AN2 AND2_1366(g8732,g8624,g7919);
  AN2 AND2_1367(g3807,g3003,g3062);
  AN2 AND2_1368(g8753,g7414,g8664);
  AN2 AND2_1369(g5848,g3860,g5519);
  AN2 AND2_1370(g8508,g8411,g7967);
  AN2 AND2_1371(g8072,g700,g7826);
  AN2 AND2_1372(g5699,g1592,g5117);
  AN2 AND2_1373(g11240,g5481,g11111);
  AN2 AND2_1374(g5398,g4610,g2224);
  AN2 AND2_1375(g6616,g6105,g3246);
  AN2 AND2_1376(g10690,g10616,g3863);
  AN2 AND2_1377(g8043,g7582,g5128);
  AN2 AND2_1378(g9590,g895,g8995);
  AN2 AND2_1379(g4128,g1976,g2779);
  AN2 AND2_1380(g6404,g2132,g5748);
  AN2 AND2_1381(g6647,g5288,g5808);
  AN2 AND2_1382(g10504,g10389,g2135);
  AN2 AND2_1383(g9657,g919,g9205);
  AN2 AND2_1384(g4542,g366,g3586);
  AN2 AND2_1385(g4330,g1163,g3693);
  AN2 AND2_1386(g3497,g2804,g1900);
  AN2 AND2_1387(g5524,g1678,g4291);
  AN2 AND2_1388(g8147,g2955,g7961);
  AN2 AND2_1389(g4554,g542,g3996);
  AN2 AND2_1390(g9899,g9889,g9367);
  AN2 AND2_1391(g5258,g700,g4756);
  AN2 AND2_1392(g7736,g6951,g3880);
  AN2 AND2_1393(g6224,g1520,g5151);
  AN2 AND2_1394(g10626,g10547,g4558);
  AN2 AND2_1395(g6320,g1292,g5949);
  AN2 AND2_1396(g7623,g664,g7079);
  AN2 AND2_1397(g10299,g8892,g10217);
  AN2 AND2_1398(g7889,g7615,g3814);
  AN2 AND2_1399(g10298,g8892,g10214);
  AN2 AND2_1400(g8413,g722,g8146);
  AN2 AND2_1401(g3979,g237,g3164);
  AN2 AND2_1402(g4902,g1848,g4243);
  AN2 AND2_1403(g5211,g1080,g4724);
  AN2 AND2_1404(g4512,g357,g3586);
  AN2 AND2_1405(g7722,g7127,g6449);
  AN2 AND2_1406(g9844,g9714,g9522);
  AN2 AND2_1407(g4490,g1141,g3913);
  AN2 AND2_1408(g4823,g207,g3946);
  AN2 AND2_1409(g6516,g5993,g3097);
  AN2 AND2_1410(g5026,g1453,g4640);
  AN2 AND2_1411(g8820,g8705,g5422);
  AN2 AND2_1412(g10737,g10687,g4840);
  AN3 AND3_45(g8936,g8115,g6778,g8849);
  AN2 AND2_1413(g10232,g8892,g10150);
  AN2 AND2_1414(g6771,g263,g5866);
  AN2 AND2_1415(g5170,g1811,g4680);
  AN2 AND2_1416(g8117,g6236,g7886);
  AN2 AND2_1417(g4529,g448,g3980);
  AN2 AND2_1418(g4348,g3497,g1909);
  AN2 AND2_1419(g9966,g9956,g9536);
  AN2 AND2_1420(g5280,g4593,g3052);
  AN2 AND2_1421(g7139,g6060,g6709);
  AN2 AND2_1422(g11099,g382,g10885);
  AN2 AND2_1423(g6892,g6472,g5805);
  AN2 AND2_1424(g9705,g1580,g9474);
  AN2 AND2_1425(g10512,g10395,g2135);
  AN2 AND2_1426(g11098,g849,g10950);
  AN2 AND2_1427(g8775,g8628,g5151);
  AN2 AND2_1428(g5083,g3709,g4586);
  AN2 AND2_1429(g5544,g1687,g4320);
  AN2 AND2_1430(g11272,g5629,g11193);
  AN2 AND2_1431(g5483,g1621,g4254);
  AN2 AND2_1432(g9948,g9928,g9392);
  AN2 AND2_1433(g4063,g2713,g2276);
  AN2 AND2_1434(g11462,g11431,g5446);
  AN2 AND2_1435(g6738,g2531,g6137);
  AN2 AND2_1436(g8060,g7593,g5919);
  AN2 AND2_1437(g6244,g2255,g5151);
  AN2 AND2_1438(g11032,g416,g10974);
  AN2 AND2_1439(g10445,g10315,g2135);
  AN2 AND2_1440(g9150,g8882,g4805);
  AN2 AND2_1441(g10316,g10223,g9097);
  AN2 AND2_1442(g5756,g1531,g5202);
  AN2 AND2_1443(g4720,g1023,g3914);
  AN2 AND2_1444(g9409,g1721,g9052);
  AN2 AND2_1445(g8995,g6454,g8929);
  AN2 AND2_1446(g6876,g4070,g6560);
  AN2 AND2_1447(g4989,g1424,g4682);
  AN2 AND2_1448(g9836,g9737,g9785);
  AN3 AND3_46(g6656,g2733,g6061,g4631);
  AN2 AND2_1449(g5514,g1941,g4284);
  AN2 AND2_1450(g8390,g8268,g6465);
  AN2 AND2_1451(g5003,g1466,g4640);
  AN2 AND2_1452(g9967,g9957,g9536);
  AN2 AND2_1453(g5145,g1639,g4673);
  AN2 AND2_1454(g4834,g219,g3946);
  AN2 AND2_1455(g4971,g1419,g4682);
  AN2 AND2_1456(g10753,g10649,g4013);
  AN2 AND2_1457(g5695,g166,g5361);
  AN2 AND2_1458(g7613,g6940,g5984);
  AN2 AND2_1459(g10736,g10658,g4840);
  AN2 AND2_1460(g11220,g962,g11054);
  AN2 AND2_1461(g7444,g7277,g5827);
  AN2 AND2_1462(g5536,g4867,g4298);
  AN2 AND2_1463(g6663,g6064,g2237);
  AN2 AND2_1464(g4670,g192,g3946);
  AN2 AND2_1465(g6824,g1371,g6596);
  AN2 AND2_1466(g4253,g1074,g3638);
  AN2 AND2_1467(g8250,g2771,g7907);
  AN2 AND2_1468(g8163,g7960,g3737);
  AN2 AND2_1469(g10764,g10643,g4840);
  AN2 AND2_1470(g5757,g1552,g5203);
  AN2 AND2_1471(g10365,g10319,g2135);
  AN2 AND2_1472(g8032,g7385,g7438);
  AN2 AND2_1473(g11591,g2988,g11561);
  AN2 AND2_1474(g8053,g7583,g5919);
  AN2 AND2_1475(g11147,g321,g10929);
  AN2 AND2_1476(g5522,g1633,g4289);
  AN2 AND2_1477(g5115,g1394,g4572);
  AN2 AND2_1478(g9837,g9697,g9751);
  AN2 AND2_1479(g9620,g2653,g9240);
  AN2 AND2_1480(g11151,g327,g10931);
  AN2 AND2_1481(g11172,g486,g11112);
  AN2 AND2_1482(g7885,g7614,g3812);
  AN2 AND2_1483(g6064,g5398,g2230);
  AN3 AND3_47(g8929,g8095,g6368,g8828);
  AN2 AND2_1484(g5595,g1621,g4524);
  AN2 AND2_1485(g5537,g4143,g4299);
  AN2 AND2_1486(g9842,g9708,g9516);
  AN2 AND2_1487(g4141,g2707,g3051);
  AN2 AND2_1488(g4341,g339,g3586);
  AN2 AND2_1489(g9192,g6454,g8955);
  AN2 AND2_1490(g7679,g1950,g6863);
  AN2 AND2_1491(g7378,g6990,g3880);
  AN2 AND2_1492(g5612,g1627,g4543);
  AN2 AND2_1493(g3939,g213,g3164);
  AN2 AND2_1494(g7135,g869,g6355);
  AN2 AND2_1495(g10970,g10852,g3390);
  AN2 AND2_1496(g11025,g426,g10974);
  AN2 AND2_1497(g9854,g9730,g9566);
  AN2 AND2_1498(g7182,g1878,g6720);
  AN2 AND2_1499(g9941,g9921,g9367);
  AN2 AND2_1500(g6194,g554,g5043);
  AN2 AND2_1501(g5128,g4474,g2733);
  AN2 AND2_1502(g4962,g1651,g4461);
  AN2 AND2_1503(g4358,g1209,g3747);
  AN2 AND2_1504(g8683,g4803,g8549);
  AN2 AND2_1505(g4506,g1113,g3944);
  AN2 AND2_1506(g6471,g5224,g6014);
  AN2 AND2_1507(g8778,g8688,g2317);
  AN2 AND2_1508(g11281,g4948,g11202);
  AN2 AND2_1509(g8735,g7600,g8632);
  AN2 AND2_1510(g11146,g318,g10928);
  AN2 AND2_1511(g3904,g2948,g2779);
  AN2 AND2_1512(g8075,g727,g7826);
  AN2 AND2_1513(g9829,g9723,g9785);
  AN3 AND3_48(g8949,g8255,g6368,g8828);
  AN2 AND2_1514(g7632,g7184,g5574);
  AN2 AND2_1515(g11290,g11246,g4226);
  AN2 AND2_1516(g6350,g5837,g4435);
  AN2 AND2_1517(g10599,g10534,g4365);
  AN2 AND2_1518(g5902,g2555,g4977);
  AN4 AND4_15(I6337,g201,g2421,g2407,g2396);
  AN2 AND2_1519(g2276,g1765,g1610);
  AN2 AND2_1520(g6438,g5853,g5797);
  AN2 AND2_1521(g5512,g1660,g4281);
  AN2 AND2_1522(g5090,g1781,g4592);
  AN2 AND2_1523(g7719,g718,g7227);
  AN2 AND2_1524(g2561,g742,g741);
  AN2 AND2_1525(g3695,g1712,g3015);
  AN2 AND2_1526(g8603,g3983,g8548);
  AN2 AND2_1527(g8039,g7587,g5128);
  AN2 AND2_1528(g9610,g925,g9192);
  AN2 AND2_1529(g3536,g2390,g3103);
  AN2 AND2_1530(g5529,g4129,g4288);
  AN2 AND2_1531(g5148,g3088,g4671);
  AN2 AND2_1532(g9124,g8881,g4802);
  AN2 AND2_1533(g9324,g8879,g5708);
  AN2 AND2_1534(g4559,g2034,g3829);
  AN2 AND2_1535(g10561,g10549,g4583);
  AN2 AND2_1536(g5698,g1571,g5116);
  AN2 AND2_1537(g11226,g461,g11057);
  AN2 AND2_1538(g10295,g8892,g10208);
  AN2 AND2_1539(g5260,g1092,g4758);
  AN2 AND2_1540(g10680,g10564,g3586);
  AN2 AND2_1541(g6822,g231,g6596);
  AN2 AND2_1542(g4905,g1853,g4243);
  AN2 AND2_1543(g11551,g11538,g4013);
  AN2 AND2_1544(g3047,g1227,g2306);
  AN2 AND2_1545(g9849,g293,g9768);
  AN2 AND2_1546(g5279,g1766,g4783);
  AN2 AND2_1547(g8404,g686,g8129);
  AN2 AND2_1548(g5720,g170,g5361);
  AN2 AND2_1549(g5318,g4401,g1857);
  AN2 AND2_1550(g8764,g7443,g8684);
  AN2 AND2_1551(g11376,g11318,g4277);
  AN2 AND2_1552(g11297,g5490,g11242);
  AN2 AND2_1553(g9898,g9887,g9367);
  OR2 OR2_0(g6895,g6776,g4875);
  OR2 OR2_1(g7189,g6632,g6053);
  OR2 OR2_2(g9510,g9125,g9111);
  OR2 OR2_3(g7297,g7132,g6323);
  OR2 OR2_4(g9088,g8927,g8381);
  OR2 OR2_5(g9923,g9865,g9707);
  OR2 OR2_6(g6485,g5848,g5067);
  OR2 OR2_7(g8771,g5483,g8652);
  OR2 OR2_8(g5813,g5617,g4869);
  OR2 OR2_9(g7963,g7687,g7182);
  OR2 OR2_10(g10643,g10624,g7736);
  OR3 OR3_0(g9886,g9607,g9592,g9759);
  OR3 OR3_1(g9951,g9902,g9899,g9803);
  OR2 OR2_11(g11625,g6535,g11597);
  OR2 OR2_12(g8945,g8801,g8710);
  OR2 OR2_13(g10489,g4961,g10367);
  OR2 OR2_14(g10559,g4141,g10512);
  OR2 OR2_15(g10558,g4126,g10510);
  OR2 OR2_16(g11338,g11283,g11178);
  OR2 OR2_17(g8435,g8403,g8075);
  OR2 OR2_18(g10544,g5511,g10495);
  OR2 OR2_19(g6911,g6342,g5681);
  OR2 OR2_20(g10865,g5538,g10752);
  OR2 OR2_21(g3698,g3121,g2480);
  OR2 OR2_22(g8214,g7472,g8004);
  OR2 OR2_23(g6124,g5181,g5188);
  OR2 OR2_24(g6469,g5698,g4959);
  OR2 OR2_25(g5587,g4714,g3904);
  OR2 OR2_26(g6177,g5444,g4712);
  OR3 OR3_2(I14585,g8995,g9205,g9192);
  OR2 OR2_27(g9891,g9741,g9760);
  OR2 OR2_28(g9913,g9849,g9691);
  OR4 OR4_0(I5600,g496,g491,g486,g481);
  OR2 OR2_29(g11257,g11234,g11019);
  OR2 OR2_30(g8236,g7526,g8001);
  OR2 OR2_31(g7385,g7235,g6746);
  OR2 OR2_32(g6898,g6790,g4881);
  OR2 OR2_33(g6900,g6787,g6246);
  OR2 OR2_34(g4264,g4048,g4053);
  OR3 OR3_3(g9726,g9411,g9420,g9489);
  OR2 OR2_35(g6088,g5260,g4522);
  OR2 OR2_36(g6923,g6353,g5695);
  OR2 OR2_37(g8194,g5168,g7940);
  OR3 OR3_4(g9676,g9454,g9292,g9274);
  OR2 OR2_38(g11256,g11186,g11018);
  OR2 OR2_39(g3860,g3107,g2167);
  OR2 OR2_40(g11280,g11254,g11153);
  OR4 OR4_1(g9727,g9650,g9663,g9362,I14866);
  OR2 OR2_41(g4997,g4581,g4584);
  OR2 OR2_42(g11624,g11595,g11571);
  OR2 OR2_43(g11300,g11213,g11091);
  OR2 OR2_44(g4238,g3999,g4007);
  OR2 OR2_45(g8814,g7945,g8728);
  OR2 OR2_46(g10401,g9317,g10291);
  OR2 OR2_47(g8773,g5491,g8653);
  OR2 OR2_48(g11231,g11156,g11013);
  OR2 OR2_49(g10864,g5532,g10751);
  OR2 OR2_50(g9624,g9316,g9313);
  OR3 OR3_5(g9953,g9945,g9939,g9669);
  OR2 OR2_51(g6122,g5172,g5180);
  OR2 OR2_52(g6465,g5825,g5041);
  OR2 OR2_53(g6934,g6363,g5720);
  OR2 OR2_54(g7664,g6855,g4084);
  OR2 OR2_55(g7246,g6465,g6003);
  OR2 OR2_56(g7203,g6640,g6058);
  OR2 OR2_57(g6096,g5268,g4542);
  OR2 OR2_58(g9747,g9173,g9509);
  OR2 OR2_59(g11314,g11224,g11102);
  OR2 OR2_60(g10733,g5227,g10674);
  OR2 OR2_61(g8921,g8827,g8748);
  OR4 OR4_2(I15054,g7853,g9782,g9624,g9785);
  OR2 OR2_62(g11269,g11196,g11031);
  OR2 OR2_63(g5555,g4389,g4397);
  OR2 OR2_64(g11268,g11194,g11030);
  OR2 OR2_65(g10485,g9317,g10376);
  OR2 OR2_66(g10555,g4103,g10504);
  OR2 OR2_67(g6481,g5722,g4972);
  OR2 OR2_68(g10712,g10662,g9531);
  OR2 OR2_69(g11335,g11279,g11175);
  OR2 OR2_70(g8249,g8018,g7710);
  OR2 OR2_71(g7638,g7265,g6488);
  OR2 OR2_72(g10567,g10514,g7378);
  OR2 OR2_73(g11487,g6662,g11464);
  OR4 OR4_3(I15210,g9839,g9964,g9852,g9882);
  OR4 OR4_4(I5805,g2102,g2099,g2096,g2088);
  OR2 OR2_74(g8941,g8796,g8706);
  OR2 OR2_75(g11443,g7130,g11407);
  OR2 OR2_76(g4231,g3991,g3998);
  OR2 OR2_77(g11278,g11253,g11150);
  OR4 OR4_5(I15039,g7853,g9809,g9624,g9785);
  OR2 OR2_78(g11286,g10670,g11209);
  OR2 OR2_79(g8431,g8387,g8071);
  OR2 OR2_80(g7133,g6616,g3067);
  OR2 OR2_81(g11306,g11216,g11095);
  OR2 OR2_82(g8252,g7988,g7679);
  OR2 OR2_83(g8812,g7939,g8724);
  OR2 OR2_84(g7846,g7722,g7241);
  OR2 OR2_85(g3875,g3275,g12);
  OR2 OR2_86(g5996,g5473,g3908);
  OR2 OR2_87(g6592,g5100,g5882);
  OR2 OR2_88(g8286,g8107,g7823);
  OR2 OR2_89(g10501,g4161,g10445);
  OR2 OR2_90(g10728,g4973,g10642);
  OR2 OR2_91(g8270,g7894,g3434);
  OR2 OR2_92(g7290,g7046,g6316);
  OR2 OR2_93(g6068,g5220,g4497);
  OR2 OR2_94(g6468,g5690,g4950);
  OR2 OR2_95(g11217,g11144,g11005);
  OR2 OR2_96(g11478,g6532,g11455);
  OR4 OR4_6(g9536,g9335,g9331,g9328,g9324);
  OR2 OR2_97(g5981,g5074,g4383);
  OR2 OR2_98(g11486,g6654,g11463);
  OR2 OR2_99(g8377,g8185,g7958);
  OR2 OR2_100(g8206,g7459,g8007);
  OR2 OR2_101(g11580,g11413,g11544);
  OR2 OR2_102(g8287,g8117,g7824);
  OR2 OR2_103(g11223,g11147,g11008);
  OR2 OR2_104(g9522,g9173,g9125);
  OR2 OR2_105(g8199,g7902,g7444);
  OR2 OR2_106(g5802,g5601,g4837);
  OR2 OR2_107(g11321,g11230,g11105);
  OR2 OR2_108(g6524,g5746,g4996);
  OR2 OR2_109(g10664,g10240,g10582);
  OR2 OR2_110(g7257,g6701,g4725);
  OR2 OR2_111(g7301,g7140,g6327);
  OR2 OR2_112(g10484,g9317,g10400);
  OR2 OR2_113(g10554,g4097,g10503);
  OR2 OR2_114(g8259,g8028,g7719);
  OR2 OR2_115(g11334,g11277,g11174);
  OR2 OR2_116(g8819,g7957,g8734);
  OR2 OR2_117(g8923,g8846,g8763);
  OR2 OR2_118(g8488,g3664,g8390);
  OR2 OR2_119(g7441,g7271,g6789);
  OR2 OR2_120(g6026,g5507,g3970);
  OR2 OR2_121(g10799,g6225,g10769);
  OR2 OR2_122(g10798,g6217,g10768);
  OR2 OR2_123(g10805,g10759,g10760);
  OR2 OR2_124(g10732,g4358,g10661);
  OR2 OR2_125(g6061,g5204,g4);
  OR2 OR2_126(g9512,g9151,g9125);
  OR2 OR2_127(g10013,I15214,I15215);
  OR2 OR2_128(g8806,g7931,g8718);
  OR2 OR2_129(g8943,g8837,g8749);
  OR2 OR2_130(g11293,g11211,g10818);
  OR2 OR2_131(g11265,g11189,g11027);
  OR2 OR2_132(g8887,g8842,g8755);
  OR2 OR2_133(g5838,g5612,g4866);
  OR2 OR2_134(g6514,g5738,g4992);
  OR2 OR2_135(g8322,g8136,g6891);
  OR2 OR2_136(g8230,g7515,g7991);
  OR2 OR2_137(g5809,g5611,g4865);
  OR2 OR2_138(g8433,g8399,g8073);
  OR2 OR2_139(g11579,g5123,g11551);
  OR2 OR2_140(g10771,g5533,g10684);
  OR2 OR2_141(g11615,g11601,g11592);
  OR2 OR2_142(g9367,g9335,g9331);
  OR3 OR3_6(g9872,g9617,g9594,g9750);
  OR2 OR2_143(g6522,g5744,g4994);
  OR2 OR2_144(g8266,g7885,g3412);
  OR2 OR2_145(g10414,g10300,g9534);
  OR2 OR2_146(g11275,g11248,g11148);
  OR2 OR2_147(g11430,g11387,g4006);
  OR2 OR2_148(g8248,g8014,g7707);
  OR3 OR3_7(g9686,g9454,g9292,g9274);
  OR2 OR2_149(g8815,g7948,g8730);
  OR2 OR2_150(g7183,g6623,g6046);
  OR2 OR2_151(g5983,g5084,g4392);
  OR2 OR2_152(g8154,g7891,g6879);
  OR2 OR2_153(g6537,g5781,g5005);
  OR2 OR2_154(g4309,g4069,g4079);
  OR2 OR2_155(g10725,g4962,g10634);
  OR2 OR2_156(g6243,g5537,g4774);
  OR4 OR4_7(I6351,g2405,g2389,g2380,g2372);
  OR3 OR3_8(g9519,g9173,g9151,g9125);
  OR2 OR2_157(g9740,g9418,g9505);
  OR2 OR2_158(g8267,g7889,g3422);
  OR3 OR3_9(g10744,g10600,g10668,I16427);
  OR2 OR2_159(g6542,g5789,g5010);
  OR2 OR2_160(g7303,g7145,g6329);
  OR2 OR2_161(g10652,g10627,g7743);
  OR2 OR2_162(g5036,g4871,g4162);
  OR2 OR2_163(g7240,g6687,g6095);
  OR2 OR2_164(g8221,g7496,g7993);
  OR2 OR2_165(g6902,g6794,g4223);
  OR3 OR3_10(I14776,g8995,g9205,g9192);
  OR2 OR2_166(g10500,g4157,g10442);
  OR2 OR2_167(g4052,g2862,g2515);
  OR4 OR4_8(I14858,g9585,g9595,g9610,g9602);
  OR2 OR2_168(g6529,g5757,g5000);
  OR2 OR2_169(g11264,g11188,g11026);
  OR4 OR4_9(I15209,g8169,g9905,g9934,g9830);
  OR2 OR2_170(g8241,g7536,g7989);
  OR2 OR2_171(g10795,g6199,g10764);
  OR2 OR2_172(g11607,g11586,g11557);
  OR2 OR2_173(g8644,g8123,g8464);
  OR3 OR3_11(g4682,g3563,g3348,g1570);
  OR2 OR2_174(g8818,g7955,g8733);
  OR2 OR2_175(g2984,g2528,g2522);
  OR2 OR2_176(g9931,g8931,g9900);
  OR2 OR2_177(g3414,g2911,g2917);
  OR2 OR2_178(g9515,g9173,g9151);
  OR2 OR2_179(g10724,g10312,g10672);
  OR2 OR2_180(g7294,g7068,g6320);
  OR2 OR2_181(g5189,g4345,g3496);
  OR2 OR2_182(g8614,g8365,g8510);
  OR2 OR2_183(g3513,g3118,g2180);
  OR2 OR2_184(g6909,g6346,g5684);
  OR4 OR4_10(I5571,g396,g391,g386,g426);
  OR2 OR2_185(g4283,g4059,g4063);
  OR2 OR2_186(g8939,g8791,g8701);
  OR2 OR2_187(g2514,I5599,I5600);
  OR2 OR2_188(g11327,g11297,g11167);
  OR2 OR2_189(g8187,g7542,g7998);
  OR2 OR2_190(g11606,g11585,g11556);
  OR2 OR2_191(g11303,g11214,g11092);
  OR2 OR2_192(g5309,g3664,g4401);
  OR3 OR3_12(g9528,g9151,g9125,g9111);
  OR2 OR2_193(g8200,g7535,g8008);
  OR3 OR3_13(g2522,g833,g829,I5629);
  OR4 OR4_11(g2315,g1163,g1166,g1113,I5363);
  OR2 OR2_194(g6506,g5731,g4989);
  OR2 OR2_195(g10649,g10626,g7741);
  OR2 OR2_196(g8159,g7895,g6886);
  OR2 OR2_197(g7626,g7060,g5267);
  OR2 OR2_198(g10770,g5525,g10682);
  OR2 OR2_199(g9566,g9052,g9030);
  OR2 OR2_200(g11483,g6633,g11460);
  OR2 OR2_201(g8811,g7935,g8722);
  OR3 OR3_14(g8642,g5236,g5205,g8465);
  OR2 OR2_202(g6545,g5795,g5025);
  OR2 OR2_203(g10767,g5500,g10681);
  OR2 OR2_204(g11326,g11296,g11166);
  OR2 OR2_205(g10898,g4220,g10777);
  OR2 OR2_206(g11252,g11099,g10969);
  OR2 OR2_207(g10719,g10303,g10666);
  OR2 OR2_208(g4609,g3400,g119);
  OR2 OR2_209(g6507,g5732,g4990);
  OR2 OR2_210(g10718,g6238,g10706);
  OR2 OR2_211(g10521,I16148,I16149);
  OR2 OR2_212(g7075,g5104,g6530);
  OR2 OR2_213(g7292,g7055,g6318);
  OR2 OR2_214(g10861,g5523,g10745);
  OR2 OR2_215(g8417,g8246,g7721);
  OR2 OR2_216(g6515,g5739,g4993);
  OR4 OR4_12(I14855,g9583,g9593,g9601,g9596);
  OR4 OR4_13(I15205,g9838,g9963,g9850,g9878);
  OR4 OR4_14(I15051,g7853,g9673,g9624,g9785);
  OR3 OR3_15(g9724,g9409,g9419,g9615);
  OR2 OR2_217(g6528,g5756,g4999);
  OR2 OR2_218(g8823,g8778,g8693);
  OR2 OR2_219(g7503,g6887,g6430);
  OR2 OR2_220(g8148,g7884,g6872);
  OR2 OR2_221(g8649,g8499,g4519);
  OR2 OR2_222(g3584,g2863,g2516);
  OR2 OR2_223(g10776,g5544,g10758);
  OR3 OR3_16(g9680,g9454,g9292,g9274);
  OR2 OR2_224(g10859,g5512,g10742);
  OR3 OR3_17(I14866,g9590,g9609,g9619);
  OR2 OR2_225(g7299,g7138,g6325);
  OR2 OR2_226(g10858,g5501,g10741);
  OR2 OR2_227(g8193,g5145,g7937);
  OR3 OR3_18(g9511,g9151,g9125,g9111);
  OR2 OR2_228(g7738,g7200,g6738);
  OR2 OR2_229(g7244,g6699,g4720);
  OR2 OR2_230(g3425,g2895,g2910);
  OR2 OR2_231(g7478,g6884,g6423);
  OR3 OR3_19(g9714,g9664,g9366,g9654);
  OR2 OR2_232(g10025,I15224,I15225);
  OR2 OR2_233(g6908,g6345,g4229);
  OR2 OR2_234(g5028,g4836,g4128);
  OR2 OR2_235(g8253,g8023,g7718);
  OR2 OR2_236(g8938,g8789,g8699);
  OR2 OR2_237(g8813,g7943,g8726);
  OR2 OR2_238(g9736,g9430,g9416);
  OR2 OR2_239(g9968,I15171,I15172);
  OR2 OR2_240(g8552,g8217,g8388);
  OR2 OR2_241(g5910,g5023,g4341);
  OR2 OR2_242(g11249,g6162,g11143);
  OR2 OR2_243(g11482,g6628,g11459);
  OR4 OR4_15(g9722,g9612,g9643,g9410,I14855);
  OR4 OR4_16(I15204,g8168,g9904,g9933,g9829);
  OR2 OR2_244(g7236,g6684,g6092);
  OR3 OR3_20(I14596,g8995,g9205,g9192);
  OR2 OR2_245(g8645,g8127,g8469);
  OR2 OR2_246(g11647,g6622,g11637);
  OR2 OR2_247(g6777,g5691,g5052);
  OR3 OR3_21(g9737,g9657,g9658,g9655);
  OR4 OR4_17(I16149,g10472,g10470,g10468,g10467);
  OR2 OR2_248(g11233,g11085,g10946);
  OR2 OR2_249(g8607,g8406,g8554);
  OR4 OR4_18(I16148,g10386,g10384,g10476,g10474);
  OR2 OR2_250(g8158,g7893,g6883);
  OR2 OR2_251(g5846,g4932,g4236);
  OR2 OR2_252(g5396,g4481,g3684);
  OR2 OR2_253(g5803,g5575,g4820);
  OR2 OR2_254(g11331,g11272,g11171);
  OR2 OR2_255(g7295,g7071,g6321);
  OR2 OR2_256(g6541,g5788,g5009);
  OR2 OR2_257(g8615,g8413,g8557);
  OR2 OR2_258(g9742,g9173,g9528);
  OR2 OR2_259(g9926,g9868,g9715);
  OR2 OR2_260(g9754,g9173,g9511);
  OR2 OR2_261(g8284,g8102,g7821);
  OR2 OR2_262(g2204,g1393,g1394);
  OR2 OR2_263(g7471,g6880,g6416);
  OR2 OR2_264(g7242,g6693,g6098);
  OR2 OR2_265(g5847,g5626,g4877);
  OR2 OR2_266(g6901,g6788,g6247);
  OR2 OR2_267(g8559,g8380,g4731);
  OR3 OR3_22(g9729,g9618,g9357,g9656);
  OR2 OR2_268(g10860,g5513,g10743);
  OR2 OR2_269(g9927,g9869,g9716);
  OR2 OR2_270(g10497,g5052,g10396);
  OR4 OR4_19(g9885,g9739,g9598,g9662,g9746);
  OR4 OR4_20(g2528,g861,g857,g853,g849);
  OR2 OR2_271(g11229,g11154,g11012);
  OR2 OR2_272(g8973,g8821,g8735);
  OR2 OR2_273(g10658,g10595,g7674);
  OR2 OR2_274(g10339,g10232,g9556);
  OR4 OR4_21(I5363,g1149,g1153,g1157,g1160);
  OR2 OR2_275(g11310,g11220,g11100);
  OR2 OR2_276(g6500,g5725,g4986);
  OR2 OR2_277(g10855,g6075,g10736);
  OR2 OR2_278(g9916,g9855,g9694);
  OR2 OR2_279(g10411,g10299,g9529);
  OR2 OR2_280(g11603,g11582,g11553);
  OR4 OR4_22(I5357,g1265,g1260,g1255,g1250);
  OR2 OR2_281(g9560,g9052,g9030);
  OR2 OR2_282(g6672,g5941,g5259);
  OR3 OR3_23(g9873,g9623,g9599,g9758);
  OR2 OR2_283(g6523,g5745,g4995);
  OR2 OR2_284(g10707,g5545,g10686);
  OR4 OR4_23(I5626,g521,g525,g530,g534);
  OR2 OR2_285(g9579,g9052,g9030);
  OR2 OR2_286(g7298,g7136,g6324);
  OR2 OR2_287(g6551,g5804,g5031);
  OR2 OR2_288(g6099,g5273,g4550);
  OR2 OR2_289(g8282,g8101,g7819);
  OR2 OR2_290(g9917,g9856,g9695);
  OR4 OR4_24(I15057,g7853,g9680,g9624,g9785);
  OR2 OR2_291(g7219,g6661,g6076);
  OR2 OR2_292(g10019,I15219,I15220);
  OR2 OR2_293(g5857,g5418,g4670);
  OR4 OR4_25(g9725,g9642,g9659,g9616,I14862);
  OR2 OR2_294(g11298,g11212,g11087);
  OR2 OR2_295(g10402,g10295,g9554);
  OR4 OR4_26(g2521,g538,g542,g476,I5626);
  OR3 OR3_24(I14751,g8995,g9205,g9192);
  OR2 OR2_296(g10866,g5539,g10753);
  OR2 OR2_297(g6534,g5772,g5003);
  OR2 OR2_298(g11232,g11158,g11015);
  OR3 OR3_25(g9706,g9644,g9386,g9591);
  OR2 OR2_299(g10001,I15204,I15205);
  OR2 OR2_300(g8776,g5510,g8655);
  OR2 OR2_301(g7225,g6666,g6079);
  OR3 OR3_26(g9888,g9648,g9608,g9757);
  OR2 OR2_302(g11261,g11238,g11023);
  OR3 OR3_27(g9956,g9948,g9942,g9815);
  OR2 OR2_303(g10923,g10778,g10715);
  OR2 OR2_304(g8264,g7879,g3389);
  OR2 OR2_305(g6513,g5737,g4991);
  OR3 OR3_28(I14835,g9621,g9645,g9588);
  OR2 OR2_306(g8641,g8120,g8463);
  OR3 OR3_29(g5361,g4316,g4093,g126);
  OR2 OR2_307(g11316,g11226,g11103);
  OR4 OR4_27(I16161,g10479,g10478,g10477,g10475);
  OR2 OR2_308(g6916,g6348,g5687);
  OR2 OR2_309(g8777,g5522,g8659);
  OR4 OR4_28(g2353,g1403,g1407,g1411,g1415);
  OR2 OR2_310(g7510,g7186,g6730);
  OR3 OR3_30(g9957,g9949,g9943,g9776);
  OR2 OR2_311(g2744,I5804,I5805);
  OR2 OR2_312(g7245,g6696,g6102);
  OR2 OR2_313(g7291,g7050,g6317);
  OR2 OR2_314(g8611,g8410,g8556);
  OR4 OR4_29(I15199,g8167,g9903,g9932,g9828);
  OR2 OR2_315(g10550,g4942,g10450);
  OR2 OR2_316(g11330,g11304,g11170);
  OR2 OR2_317(g10721,g10306,g10669);
  OR2 OR2_318(g8153,g7888,g6875);
  OR2 OR2_319(g10773,g5540,g10685);
  OR2 OR2_320(g3688,g3144,g2454);
  OR4 OR4_30(I15225,g9842,g9967,g9859,g9881);
  OR2 OR2_321(g6042,g5535,g3987);
  OR2 OR2_322(g10655,g10561,g7389);
  OR2 OR2_323(g11259,g11236,g11021);
  OR2 OR2_324(g11225,g11149,g11009);
  OR2 OR2_325(g5914,g5029,g4343);
  OR2 OR2_326(g11258,g11235,g11020);
  OR2 OR2_327(g6054,g5199,g4483);
  OR3 OR3_31(g9728,g9412,g9422,g9426);
  OR3 OR3_32(g9730,g9414,g9425,g9423);
  OR2 OR2_328(g5820,g5595,g4834);
  OR3 OR3_33(g8574,g5679,g7853,g8465);
  OR2 OR2_329(g11602,g11581,g11552);
  OR2 OR2_330(g10502,g4169,g10365);
  OR2 OR2_331(g10557,g4123,g10508);
  OR4 OR4_31(I15171,g8175,g9909,g9896,g9835);
  OR2 OR2_332(g11337,g11282,g11177);
  OR2 OR2_333(g7465,g6876,g6410);
  OR2 OR2_334(g8262,g7970,g7625);
  OR2 OR2_335(g8889,g8844,g8756);
  OR2 OR2_336(g7096,g6544,g5911);
  OR2 OR2_337(g5995,g5097,g5099);
  OR2 OR2_338(g8285,g8104,g7822);
  OR2 OR2_339(g10791,g6186,g10762);
  OR2 OR2_340(g2499,I5570,I5571);
  OR3 OR3_34(I14607,g8995,g9205,g9192);
  OR2 OR2_341(g6049,g5254,g3718);
  OR2 OR2_342(g9920,g9860,g9701);
  OR2 OR2_343(g10556,g4115,g10506);
  OR2 OR2_344(g8643,g8364,g8508);
  OR2 OR2_345(g5810,g5588,g4823);
  OR2 OR2_346(g11336,g11281,g11176);
  OR2 OR2_347(g8742,g8135,g8598);
  OR2 OR2_348(g8926,g8848,g8764);
  OR2 OR2_349(g7218,g6655,g6070);
  OR4 OR4_32(I15224,g8174,g9908,g9937,g9834);
  OR2 OR2_350(g7293,g7063,g6319);
  OR2 OR2_351(g11288,g11204,g11070);
  OR2 OR2_352(g10800,g6245,g10772);
  OR2 OR2_353(g11308,g11218,g11098);
  OR2 OR2_354(g8269,g7892,g3429);
  OR2 OR2_355(g10417,g10301,g9527);
  OR2 OR2_356(g10936,g5170,g10808);
  OR2 OR2_357(g9388,g9240,g9223);
  OR2 OR2_358(g6185,g5470,g4715);
  OR2 OR2_359(g6470,g5699,g4960);
  OR2 OR2_360(g6897,g6771,g6240);
  OR2 OR2_361(g8885,g8841,g8754);
  OR2 OR2_362(g11260,g11237,g11022);
  OR2 OR2_363(g11488,g6671,g11465);
  OR2 OR2_364(g6105,g5279,g4559);
  OR2 OR2_365(g10807,g10701,g10761);
  OR2 OR2_366(g10639,g10623,g7734);
  OR2 OR2_367(g4556,g3536,g2916);
  OR2 OR2_368(g8288,g8119,g7825);
  OR2 OR2_369(g6755,g6106,g5479);
  OR3 OR3_35(I14862,g9587,g9600,g9611);
  OR4 OR4_33(I16160,g10394,g10392,g10482,g10481);
  OR4 OR4_34(I15042,g7853,g9686,g9624,g9785);
  OR2 OR2_370(g11610,g11589,g11560);
  OR4 OR4_35(g9711,g9660,g9390,g9359,g9589);
  OR2 OR2_371(g6045,g5541,g3989);
  OR2 OR2_372(g11270,g11198,g11032);
  OR2 OR2_373(g7258,g6549,g5913);
  OR2 OR2_374(g6059,g5211,g4489);
  OR2 OR2_375(g10007,I15209,I15210);
  OR2 OR2_376(g11267,g11192,g11029);
  OR2 OR2_377(g11294,g6576,g11210);
  OR3 OR3_36(g9509,g9151,g9125,g9111);
  OR2 OR2_378(g7211,g6647,g6067);
  OR2 OR2_379(g5404,g4487,g3696);
  OR2 OR2_380(g4089,g1959,g3318);
  OR4 OR4_36(I15219,g8172,g9907,g9936,g9833);
  OR2 OR2_381(g11219,g11145,g11006);
  OR2 OR2_382(g6015,g5497,g3942);
  OR2 OR2_383(g10720,g10304,g10667);
  OR2 OR2_384(g8265,g7881,g3396);
  OR2 OR2_385(g5224,g4360,g3512);
  OR3 OR3_37(g9700,g9358,g9667,I14827);
  OR2 OR2_386(g7106,g6554,g5917);
  OR2 OR2_387(g8770,g5476,g8651);
  OR2 OR2_388(g11201,g11152,g11011);
  OR3 OR3_38(g9950,g9901,g9898,g9779);
  OR4 OR4_37(g9723,g9620,g9652,g9391,I14858);
  OR2 OR2_389(g2309,I5357,I5358);
  OR2 OR2_390(g11266,g11190,g11028);
  OR2 OR2_391(g10727,g4969,g10638);
  OR2 OR2_392(g10863,g5531,g10750);
  OR2 OR2_393(g8429,g8385,g8069);
  OR2 OR2_394(g9751,g9515,g9510);
  OR2 OR2_395(g8281,g8097,g7818);
  OR2 OR2_396(g6910,g6341,g5680);
  OR2 OR2_397(g8639,g8118,g8462);
  OR3 OR3_39(g9673,g9454,g9292,g9274);
  OR2 OR2_398(g11285,g11255,g11161);
  OR2 OR2_399(g11305,g11215,g11093);
  OR4 OR4_38(I15177,g9844,g9960,g9863,g9876);
  OR3 OR3_40(g9734,g9415,g9428,g9421);
  OR3 OR3_41(I14827,g9603,g9614,g9584);
  OR2 OR2_400(g5824,g5602,g4839);
  OR2 OR2_401(g8715,g8416,g8687);
  OR2 OR2_402(g5762,g5178,g5186);
  OR2 OR2_403(g6538,g5782,g5006);
  OR2 OR2_404(g5590,g4718,g4723);
  OR2 OR2_405(g10726,g10316,g10673);
  OR2 OR2_406(g3120,I6350,I6351);
  OR2 OR2_407(g9573,g9052,g9030);
  OR3 OR3_42(g4640,g3348,g3563,g1527);
  OR2 OR2_408(g6093,g5264,g4534);
  OR2 OR2_409(g8162,g7898,g6889);
  OR2 OR2_410(g8268,g7962,g7613);
  OR2 OR2_411(g9569,g9052,g9030);
  OR2 OR2_412(g11485,g6646,g11462);
  OR2 OR2_413(g10797,g6206,g10766);
  OR3 OR3_43(I14779,g8995,g9205,g9192);
  OR2 OR2_414(g10408,g10298,g9553);
  OR2 OR2_415(g10635,g10622,g7732);
  OR2 OR2_416(g2305,I5351,I5352);
  OR4 OR4_39(I15176,g8176,g9910,g9897,g9836);
  OR2 OR2_417(g3435,g2945,g2950);
  OR2 OR2_418(g9924,g9866,g9709);
  OR2 OR2_419(g10711,g5547,g10690);
  OR2 OR2_420(g5814,g5591,g4827);
  OR2 OR2_421(g5038,g4878,g4884);
  OR4 OR4_40(I15215,g9840,g9965,g9854,g9879);
  OR2 OR2_422(g8226,g7504,g8002);
  OR2 OR2_423(g7367,g7224,g6744);
  OR2 OR2_424(g7457,g6873,g6404);
  OR2 OR2_425(g5229,g4364,g3516);
  OR2 OR2_426(g5993,g5090,g4400);
  OR2 OR2_427(g8283,g8098,g7820);
  OR2 OR2_428(g7971,g5110,g7549);
  OR2 OR2_429(g8602,g8401,g8550);
  OR2 OR2_430(g8920,g8845,g8759);
  OR2 OR2_431(g10663,g10237,g10581);
  OR2 OR2_432(g6074,g5349,g1);
  OR2 OR2_433(g8261,g7876,g3383);
  OR2 OR2_434(g10862,g5524,g10746);
  OR2 OR2_435(g5837,g5640,g4224);
  OR2 OR2_436(g11333,g11274,g11173);
  OR2 OR2_437(g6080,g5249,g4512);
  OR2 OR2_438(g6480,g5721,g4971);
  OR2 OR2_439(g7740,g7209,g6741);
  OR2 OR2_440(g10702,g10562,g3877);
  OR3 OR3_44(g9697,g9665,g9606,I14822);
  OR2 OR2_441(g8203,g7453,g7999);
  OR2 OR2_442(g9914,g9851,g9692);
  OR2 OR2_443(g10564,g10560,g7368);
  OR2 OR2_444(g11484,g6639,g11461);
  OR2 OR2_445(g5842,g5618,g4870);
  OR4 OR4_41(I15200,g9837,g9962,g9848,g9880);
  OR2 OR2_446(g11609,g11588,g11559);
  OR3 OR3_45(I14582,g8995,g9205,g9192);
  OR2 OR2_447(g8940,g8793,g8703);
  OR2 OR2_448(g11312,g11222,g11101);
  OR2 OR2_449(g11608,g11587,g11558);
  OR2 OR2_450(g6000,g5480,g3912);
  OR2 OR2_451(g8428,g8382,g8068);
  OR2 OR2_452(g8430,g8386,g8070);
  OR2 OR2_453(g9922,g9864,g9705);
  OR2 OR2_454(g8247,g8010,g7704);
  OR2 OR2_455(g3438,g2939,g2944);
  OR4 OR4_42(I5576,g431,g435,g440,g444);
  OR2 OR2_456(g6924,g6362,g4261);
  OR2 OR2_457(g5405,g4476,g3440);
  OR2 OR2_458(g8638,g8108,g8461);
  OR2 OR2_459(g8609,g8408,g8555);
  OR2 OR2_460(g9995,I15199,I15200);
  OR2 OR2_461(g8883,g8838,g8753);
  OR4 OR4_43(I15214,g8170,g9906,g9935,g9831);
  OR3 OR3_46(g2538,g1466,g1458,I5649);
  OR2 OR2_462(g11329,g11302,g11169);
  OR2 OR2_463(g4255,g4009,g4047);
  OR2 OR2_464(g11328,g11299,g11168);
  OR3 OR3_47(g9704,g9385,g9605,I14835);
  OR4 OR4_44(I5352,g1129,g1125,g1121,g1117);
  OR2 OR2_465(g8774,g5499,g8654);
  OR3 OR3_48(g9954,g9946,g9940,g9781);
  OR2 OR2_466(g10405,g10297,g9530);
  OR2 OR2_467(g9363,g9205,g9192);
  OR2 OR2_468(g5849,g4949,g4260);
  OR4 OR4_45(I5599,g516,g511,g506,g501);
  OR2 OR2_469(g7204,g6645,g6062);
  OR2 OR2_470(g7300,g7139,g6326);
  OR2 OR2_471(g4293,g4064,g4068);
  OR2 OR2_472(g9912,g9847,g9690);
  OR2 OR2_473(g6533,g5771,g5002);
  OR2 OR2_474(g8816,g7951,g8731);
  OR2 OR2_475(g9929,g9871,g9718);
  OR2 OR2_476(g5819,g5625,g4876);
  OR3 OR3_49(I14831,g9613,g9622,g9586);
  OR2 OR2_477(g5852,g5632,g4883);
  OR2 OR2_478(g8263,g8032,g7720);
  OR2 OR2_479(g3431,g2951,g2957);
  OR3 OR3_50(g9683,g9454,g9292,g9274);
  OR2 OR2_480(g8631,g8474,g7449);
  OR2 OR2_481(g6922,g6352,g5694);
  OR2 OR2_482(g8817,g7954,g8732);
  OR4 OR4_46(g9735,g9649,g9651,g9384,g9361);
  OR2 OR2_483(g8605,g8404,g8553);
  OR2 OR2_484(g11263,g11187,g11025);
  OR2 OR2_485(g6739,g5769,g5780);
  OR2 OR2_486(g11332,g11273,g11172);
  OR2 OR2_487(g7143,g6619,g6039);
  OR2 OR2_488(g6479,g5707,g4968);
  OR4 OR4_47(I15048,g7853,g9683,g9624,g9785);
  OR2 OR2_489(g6501,g5726,g4987);
  OR3 OR3_51(g9702,g9365,g9647,I14831);
  OR2 OR2_490(g11221,g11146,g11007);
  OR3 OR3_52(g9952,g9944,g9938,g9817);
  OR2 OR2_491(g11613,g11600,g11591);
  OR2 OR2_492(g7621,g5108,g6994);
  OR2 OR2_493(g3399,g2918,g2940);
  OR2 OR2_494(g11605,g11584,g11555);
  OR2 OR2_495(g4274,g4054,g4058);
  OR3 OR3_53(I14602,g8995,g9205,g9192);
  OR4 OR4_48(I15033,g7853,g9804,g9624,g9785);
  OR2 OR2_496(g10717,g6235,g10705);
  OR3 OR3_54(I5629,g845,g841,g837);
  OR2 OR2_497(g9925,g9867,g9712);
  OR2 OR2_498(g3819,g3275,g9);
  OR2 OR2_499(g6912,g6350,g4235);
  OR2 OR2_500(g10723,g4952,g10633);
  OR2 OR2_501(g6929,g6360,g5704);
  OR2 OR2_502(g10646,g10625,g7739);
  OR2 OR2_503(g9516,g9151,g9125);
  OR2 OR2_504(g6626,g5934,g123);
  OR4 OR4_49(I6350,g2445,g2437,g2433,g2419);
  OR2 OR2_505(g11325,g11295,g11165);
  OR4 OR4_50(I5366,g1280,g1284,g1292,g1296);
  OR3 OR3_55(I5649,g1499,g1486,g1482);
  OR2 OR2_506(g6894,g6763,g4868);
  OR3 OR3_56(g9738,g9417,g9447,g9506);
  OR2 OR2_507(g8383,g8163,g5051);
  OR2 OR2_508(g8779,g5530,g8663);
  OR2 OR2_509(g8161,g8005,g7185);
  OR2 OR2_510(g8451,g3440,g8366);
  OR2 OR2_511(g9915,g9853,g9693);
  OR4 OR4_51(g2316,g1300,g1304,g1270,I5366);
  OR2 OR2_512(g5576,g4675,g3664);
  OR2 OR2_513(g10857,g6090,g10738);
  OR2 OR2_514(g10793,g6194,g10763);
  OR2 OR2_515(g7511,g6890,g6438);
  OR2 OR2_516(g8944,g8799,g8708);
  OR2 OR2_517(g10765,g5492,g10680);
  OR2 OR2_518(g10549,g4951,g10451);
  OR2 OR2_519(g7092,g6540,g5902);
  OR2 OR2_520(g11604,g11583,g11554);
  OR2 OR2_521(g8434,g8400,g8074);
  OR2 OR2_522(g6546,g5796,g5026);
  OR2 OR2_523(g3354,g2920,g2124);
  OR2 OR2_524(g9928,g9870,g9717);
  OR2 OR2_525(g11262,g11240,g11024);
  OR4 OR4_52(g9785,g9010,g8995,g9388,g9363);
  OR2 OR2_526(g5867,g3440,g4921);
  OR2 OR2_527(g8210,g7466,g7995);
  OR2 OR2_528(g10533,g4933,g10449);
  OR2 OR2_529(g9563,g9052,g9030);
  OR2 OR2_530(g6906,g6791,g5674);
  OR2 OR2_531(g7375,g7230,g6745);
  OR2 OR2_532(g7651,g7135,g4084);
  OR4 OR4_53(I5570,g416,g411,g406,g401);
  OR3 OR3_57(g9731,g9641,g9364,g9387);
  OR2 OR2_533(g11247,g11097,g10949);
  OR4 OR4_54(I15045,g7853,g9676,g9624,g9785);
  OR2 OR2_534(g10856,g6083,g10737);
  OR2 OR2_535(g9557,g9052,g9030);
  OR2 OR2_536(g7184,g6625,g6047);
  OR2 OR2_537(g11612,g11599,g11590);
  OR2 OR2_538(g7384,g7088,g6618);
  OR2 OR2_539(g11324,g11271,g11164);
  OR2 OR2_540(g8922,g8822,g8736);
  OR4 OR4_55(I5358,g1245,g1240,g1235,g1275);
  OR3 OR3_58(g9955,g9947,g9941,g9808);
  OR4 OR4_56(g2501,g448,g452,g421,I5576);
  OR2 OR2_541(g7231,g6673,g6087);
  OR2 OR2_542(g6078,g4503,g5256);
  OR2 OR2_543(g6478,g5706,g4967);
  OR2 OR2_544(g6907,g6792,g5675);
  OR2 OR2_545(g6035,g5518,g3974);
  OR2 OR2_546(g8937,g8786,g8698);
  OR2 OR2_547(g7742,g7217,g6743);
  OR2 OR2_548(g10722,g10308,g10671);
  OR2 OR2_549(g9918,g9858,g9698);
  OR2 OR2_550(g5403,g4486,g3695);
  OR2 OR2_551(g7926,g7435,g6892);
  OR2 OR2_552(g6915,g6347,g5686);
  OR2 OR2_553(g5841,g4914,g4230);
  OR4 OR4_57(I15220,g9841,g9966,g9857,g9877);
  OR2 OR2_554(g10529,I16160,I16161);
  OR2 OR2_555(g11246,g11094,g10948);
  OR2 OR2_556(g6002,g5489,g3939);
  OR2 OR2_557(g7712,g7125,g3540);
  OR2 OR2_558(g8810,g7933,g8720);
  OR2 OR2_559(g9921,g9862,g9703);
  OR2 OR2_560(g8432,g8389,g8072);
  OR4 OR4_58(I15172,g9843,g9959,g9861,g9874);
  OR3 OR3_59(I14822,g9597,g9604,g9582);
  OR2 OR2_561(g6928,g6359,g5703);
  OR2 OR2_562(g8157,g7965,g7623);
  OR2 OR2_563(g6930,g6364,g4269);
  OR2 OR2_564(g7660,g7059,g6583);
  OR2 OR2_565(g6899,g6463,g5471);
  OR2 OR2_566(g9392,g9328,g9324);
  OR2 OR2_567(g11318,g11228,g11104);
  OR3 OR3_60(I16427,g10683,g10608,g10604);
  OR2 OR2_568(g11227,g11151,g11010);
  OR2 OR2_569(g11058,g10933,g5280);
  OR4 OR4_59(I5351,g1145,g1141,g1137,g1133);
  OR3 OR3_61(g9708,g9653,g9389,g9646);
  OR2 OR2_570(g6071,g5228,g4505);
  OR2 OR2_571(g9911,g9846,g9689);
  OR2 OR2_572(g7102,g6550,g5915);
  OR2 OR2_573(g7302,g7141,g6328);
  OR2 OR2_574(g6038,g5528,g3979);
  OR2 OR2_575(g4239,g4000,g4008);
  OR2 OR2_576(g8646,g8224,g8547);
  OR2 OR2_577(g9974,I15176,I15177);
  OR2 OR2_578(g5823,g5631,g4882);
  OR2 OR2_579(g6918,g6358,g4252);
  OR2 OR2_580(g7265,g6756,g6204);
  OR4 OR4_60(I5804,g2111,g2109,g2106,g2104);
  OR2 OR2_581(g5851,g4941,g4253);
  OR2 OR2_582(g11481,g6624,g11458);
  OR2 OR2_583(g10336,g10230,g9572);
  OR2 OR2_584(g7296,g7131,g6322);
  OR2 OR2_585(g4300,g3546,g2391);
  OR2 OR2_586(g8647,g8130,g8470);
  ND2 NAND2_0(g8546,g3983,g8390);
  ND2 NAND2_1(g2516,I5612,I5613);
  ND2 NAND2_2(g2987,g2481,g883);
  ND2 NAND2_3(I5593,g1703,I5591);
  ND2 NAND2_4(g8970,g5548,g8839);
  ND2 NAND2_5(I10519,g6231,g822);
  ND2 NAND2_6(I11279,g305,I11278);
  ND4 NAND4_0(g7990,g7011,g6995,g7562,g7550);
  ND2 NAND2_7(I11278,g305,g6485);
  ND2 NAND2_8(g3978,g3207,g1822);
  ND2 NAND2_9(I5264,g456,I5263);
  ND2 NAND2_10(I8640,g4278,g516);
  ND2 NAND2_11(I6761,g2943,I6760);
  ND2 NAND2_12(I17400,g11418,g11416);
  ND2 NAND2_13(I5450,g1235,I5449);
  ND2 NAND2_14(I16060,g10372,I16058);
  ND2 NAND2_15(I6746,g2938,g1453);
  ND2 NAND2_16(I11975,g1462,I11973);
  ND2 NAND2_17(I12136,g7110,g131);
  ND2 NAND2_18(I11937,g1458,I11935);
  ND2 NAND2_19(g2959,I6167,I6168);
  ND2 NAND2_20(I5878,g2120,g2115);
  ND2 NAND2_21(g2517,I5619,I5620);
  ND2 NAND2_22(g5552,g4777,g4401);
  ND2 NAND2_23(I6468,g23,I6467);
  ND2 NAND2_24(I8796,g4672,I8795);
  ND2 NAND2_25(g10392,I15891,I15892);
  ND2 NAND2_26(I5611,g1280,g1284);
  ND2 NAND2_27(g8738,g8688,g4921);
  ND2 NAND2_28(I6716,g201,I6714);
  ND2 NAND2_29(g2310,g591,g605);
  ND2 NAND2_30(I7685,g3460,I7683);
  ND2 NAND2_31(g3056,g2374,g599);
  ND2 NAND2_32(I12108,g135,I12106);
  ND3 NAND3_0(g3529,g2310,g3062,g2325);
  ND2 NAND2_33(I6747,g2938,I6746);
  ND2 NAND2_34(g2236,I5230,I5231);
  ND2 NAND2_35(g7584,I12075,I12076);
  ND2 NAND2_36(I15870,g10358,g2713);
  ND2 NAND2_37(I16067,g2765,I16065);
  ND2 NAND2_38(I7562,g3533,g654);
  ND2 NAND2_39(I13531,g8253,I13529);
  ND2 NAND2_40(I8797,g1145,I8795);
  ND2 NAND2_41(I17584,g11354,g11515);
  ND2 NAND2_42(I11936,g7004,I11935);
  ND2 NAND2_43(I15257,g9984,I15256);
  ND2 NAND2_44(g8402,I13505,I13506);
  ND3 NAND3_1(g8824,g8502,g8501,g8739);
  ND2 NAND2_45(I6186,g2511,g466);
  ND2 NAND2_46(g11496,I17504,I17505);
  ND2 NAND2_47(I16001,g2683,I15999);
  ND2 NAND2_48(I6125,g2215,I6124);
  ND2 NAND2_49(I11909,g1474,I11907);
  ND2 NAND2_50(I12040,g1466,I12038);
  ND2 NAND2_51(I13909,g1432,I13907);
  ND2 NAND2_52(g3625,I6771,I6772);
  ND2 NAND2_53(I11908,g6967,I11907);
  ND2 NAND2_54(g10470,I16008,I16009);
  ND2 NAND2_55(I13908,g8526,I13907);
  ND2 NAND2_56(g3813,I7034,I7035);
  ND2 NAND2_57(I8650,g4824,g778);
  ND2 NAND2_58(g6207,I9947,I9948);
  ND2 NAND2_59(I16066,g10428,I16065);
  ND2 NAND2_60(g2948,I6144,I6145);
  ND2 NAND2_61(I11242,g6760,I11241);
  ND2 NAND2_62(g10467,I15993,I15994);
  ND2 NAND2_63(I6187,g2511,I6186);
  ND2 NAND2_64(g6488,g6027,g6019);
  ND2 NAND2_65(I5500,g1255,g1007);
  ND2 NAND2_66(I11974,g7001,I11973);
  ND2 NAND2_67(I12062,g1478,I12060);
  ND2 NAND2_68(g5300,I8771,I8772);
  ND2 NAND2_69(I5184,g1415,g1515);
  ND2 NAND2_70(I13293,g1882,g8161);
  ND2 NAND2_71(I6200,g2525,I6199);
  ND2 NAND2_72(I13265,g1909,g8154);
  ND2 NAND2_73(I5024,g995,I5023);
  ND2 NAND2_74(I7863,g4099,g774);
  ND2 NAND2_75(g8705,I13991,I13992);
  ND2 NAND2_76(g8471,I13660,I13661);
  ND2 NAND2_77(I15256,g9984,g9980);
  ND2 NAND2_78(I6145,g646,I6143);
  ND2 NAND2_79(I13992,g8688,I13990);
  ND2 NAND2_80(I11510,g1806,I11508);
  ND2 NAND2_81(g10853,g10731,g5034);
  ND2 NAND2_82(I5231,g148,I5229);
  ND2 NAND2_83(I12047,g1486,I12045);
  ND2 NAND2_84(I10771,g1801,I10769);
  ND2 NAND2_85(g10477,I16045,I16046);
  ND2 NAND2_86(g7582,I12061,I12062);
  ND2 NAND2_87(I5104,g431,g435);
  ND2 NAND2_88(g8409,I13530,I13531);
  ND2 NAND2_89(I6447,g2264,g1776);
  ND2 NAND2_90(I4956,g327,I4954);
  ND2 NAND2_91(I5613,g1284,I5611);
  ND2 NAND2_92(I8481,g3530,I8479);
  ND2 NAND2_93(g5278,I8739,I8740);
  ND2 NAND2_94(I6880,g3301,I6879);
  ND2 NAND2_95(I15431,g10047,I15430);
  ND2 NAND2_96(g5548,g1840,g4401);
  ND4 NAND4_1(g7671,g7011,g6995,g6984,g6974);
  ND2 NAND2_97(I12020,g7119,I12019);
  ND2 NAND2_98(g10665,I16331,I16332);
  ND2 NAND2_99(I16469,g10518,I16467);
  ND2 NAND2_100(I5014,g1007,I5013);
  ND2 NAND2_101(I13523,g8249,I13521);
  ND2 NAND2_102(I16039,g2707,I16037);
  ND2 NAND2_103(I16468,g10716,I16467);
  ND2 NAND2_104(I12046,g6951,I12045);
  ND2 NAND2_105(g4476,g3807,g3071);
  ND2 NAND2_106(g10476,I16038,I16039);
  ND2 NAND2_107(I16038,g10427,I16037);
  ND2 NAND2_108(I8676,g4374,g1027);
  ND2 NAND2_109(I12113,g7093,g162);
  ND2 NAND2_110(I8761,g4616,g1129);
  ND2 NAND2_111(g3204,g2571,g2061);
  ND2 NAND2_112(I15993,g10422,I15992);
  ND2 NAND2_113(I5036,g1019,I5034);
  ND2 NAND2_114(I14263,g8843,g1814);
  ND2 NAND2_115(g8298,I13249,I13250);
  ND2 NAND2_116(I5135,g521,g525);
  ND2 NAND2_117(g2405,I5485,I5486);
  ND2 NAND2_118(I7034,g3089,I7033);
  ND2 NAND2_119(I15443,g10122,I15441);
  ND2 NAND2_120(I6166,g2236,g153);
  ND2 NAND2_121(I8624,g4267,g511);
  ND2 NAND2_122(I16015,g10425,g2695);
  ND2 NAND2_123(I8677,g4374,I8676);
  ND2 NAND2_124(I8576,g4234,I8575);
  ND2 NAND2_125(I14613,g9204,I14612);
  ND2 NAND2_126(I8716,g4601,I8715);
  ND2 NAND2_127(g3530,I6715,I6716);
  ND2 NAND2_128(g8405,I13514,I13515);
  ND4 NAND4_2(g4104,g3215,g3247,g2439,g3200);
  ND2 NAND2_129(I12003,g7082,I12002);
  ND2 NAND2_130(g2177,I5127,I5128);
  ND2 NAND2_131(g3010,g2382,g2399);
  ND2 NAND2_132(g5179,I8576,I8577);
  ND2 NAND2_133(I17395,g11414,I17393);
  ND2 NAND2_134(g7067,I11279,I11280);
  ND4 NAND4_3(g7994,g7011,g7574,g6984,g7550);
  ND2 NAND2_135(I6167,g2236,I6166);
  ND2 NAND2_136(I5265,g461,I5263);
  ND2 NAND2_137(I6989,g2760,I6988);
  ND2 NAND2_138(I13274,g8158,I13272);
  ND2 NAND2_139(I10507,g6221,g786);
  ND2 NAND2_140(I13530,g704,I13529);
  ND2 NAND2_141(I5164,g1508,g1499);
  ND2 NAND2_142(g9107,I14443,I14444);
  ND2 NAND2_143(I9559,g782,I9557);
  ND2 NAND2_144(I8577,g496,I8575);
  ND2 NAND2_145(g2510,I5592,I5593);
  ND2 NAND2_146(g8177,I13077,I13078);
  ND2 NAND2_147(I8717,g4052,I8715);
  ND2 NAND2_148(I5296,g794,I5295);
  ND2 NAND2_149(g5209,I8625,I8626);
  ND4 NAND4_4(g7950,g7395,g7390,g7380,g7273);
  ND2 NAND2_150(g2088,I4911,I4912);
  ND2 NAND2_151(I16000,g10423,I15999);
  ND2 NAND2_152(I5371,g971,g976);
  ND2 NAND2_153(g2215,I5185,I5186);
  ND2 NAND2_154(g7101,g6617,g2364);
  ND2 NAND2_155(I5675,g1218,g1223);
  ND2 NAND2_156(I8544,g4218,I8543);
  ND2 NAND2_157(g6577,I10520,I10521);
  ND2 NAND2_158(I5297,g798,I5295);
  ND2 NAND2_159(I13537,g658,g8157);
  ND2 NAND2_160(I13283,g1927,g8159);
  ND2 NAND2_161(g4749,g3710,g2061);
  ND2 NAND2_162(I11982,g1482,I11980);
  ND2 NAND2_163(I8514,g4873,I8513);
  ND2 NAND2_164(I13091,g1840,I13089);
  ND2 NAND2_165(g2943,I6125,I6126);
  ND2 NAND2_166(I15908,g10302,I15906);
  ND2 NAND2_167(I6879,g3301,g1351);
  ND2 NAND2_168(I8763,g1129,I8761);
  ND2 NAND2_169(I5449,g1235,g991);
  ND3 NAND3_2(g8825,g8502,g8738,g8506);
  ND2 NAND2_170(I16007,g10424,g2689);
  ND2 NAND2_171(I5865,g2107,g2105);
  ND2 NAND2_172(I5604,g1149,g1153);
  ND2 NAND2_173(g2433,I5517,I5518);
  ND2 NAND2_174(I6111,g1494,I6109);
  ND2 NAND2_175(g2096,I4929,I4930);
  ND2 NAND2_176(I13522,g695,I13521);
  ND2 NAND2_177(I10770,g5944,I10769);
  ND2 NAND2_178(g6027,g4566,g4921);
  ND4 NAND4_5(g7992,g7011,g7574,g6984,g6974);
  ND2 NAND2_179(I5539,g1270,I5538);
  ND2 NAND2_180(I17394,g11415,I17393);
  ND2 NAND2_181(I13553,g668,I13552);
  ND2 NAND2_182(I8642,g516,I8640);
  ND2 NAND2_183(g7573,I12046,I12047);
  ND2 NAND2_184(g11416,I17296,I17297);
  ND2 NAND2_185(g6003,g5552,g5548);
  ND2 NAND2_186(g8934,I14278,I14279);
  ND2 NAND2_187(I15992,g10422,g2677);
  ND2 NAND2_188(I7683,g1023,g3460);
  ND2 NAND2_189(I4910,g386,g318);
  ND4 NAND4_6(g3209,g2550,g2061,g2564,g2571);
  ND2 NAND2_190(I6794,g143,I6792);
  ND2 NAND2_191(I10521,g822,I10519);
  ND2 NAND2_192(I5486,g1011,I5484);
  ND2 NAND2_193(I15442,g10035,I15441);
  ND2 NAND2_194(g6858,I10931,I10932);
  ND2 NAND2_195(I5185,g1415,I5184);
  ND2 NAND2_196(g5304,I8779,I8780);
  ND2 NAND2_197(g2354,g1515,g1520);
  ND2 NAND2_198(I15615,g10043,g10153);
  ND2 NAND2_199(I17281,g11360,g11357);
  ND2 NAND2_200(I5470,g999,I5468);
  ND2 NAND2_201(I11509,g6580,I11508);
  ND2 NAND2_202(I5025,g1275,I5023);
  ND2 NAND2_203(I11508,g6580,g1806);
  ND2 NAND2_204(I15430,g10047,g10044);
  ND2 NAND2_205(I14612,g9204,g611);
  ND2 NAND2_206(g4675,g4073,g3247);
  ND2 NAND2_207(I14272,g1822,I14270);
  ND2 NAND2_208(g2979,I6208,I6209);
  ND2 NAND2_209(I17290,g11363,I17288);
  ND2 NAND2_210(g5269,I8716,I8717);
  ND2 NAND2_211(g4297,I7563,I7564);
  ND2 NAND2_212(I12002,g7082,g153);
  ND2 NAND2_213(I5006,g421,I5005);
  ND2 NAND2_214(I12128,g170,I12126);
  ND2 NAND2_215(I5105,g431,I5104);
  ND2 NAND2_216(I6323,g2050,I6322);
  ND2 NAND2_217(g7588,I12093,I12094);
  ND2 NAND2_218(I6666,g2776,I6664);
  ND2 NAND2_219(g3623,I6761,I6762);
  ND2 NAND2_220(I5373,g976,I5371);
  ND2 NAND2_221(I8529,g481,I8527);
  ND2 NAND2_222(I5283,g758,I5282);
  ND2 NAND2_223(I7224,g2981,I7223);
  ND2 NAND2_224(I5007,g312,I5005);
  ND2 NAND2_225(I5459,g1240,g1003);
  ND2 NAND2_226(I17297,g11369,I17295);
  ND3 NAND3_3(g8746,g8617,g6517,g6509);
  ND2 NAND2_227(I6143,g1976,g646);
  ND2 NAND2_228(I5015,g1011,I5013);
  ND2 NAND2_229(g8932,I14264,I14265);
  ND2 NAND2_230(I16073,g845,I16072);
  ND2 NAND2_231(I6988,g2760,g986);
  ND2 NAND2_232(g3205,g1814,g2571);
  ND2 NAND2_233(I8652,g778,I8650);
  ND2 NAND2_234(I9558,g5598,I9557);
  ND2 NAND2_235(I5203,g369,I5202);
  ND2 NAND2_236(g7533,I11936,I11937);
  ND2 NAND2_237(g3634,I6806,I6807);
  ND2 NAND2_238(I6792,g2959,g143);
  ND2 NAND2_239(g3304,I6468,I6469);
  ND2 NAND2_240(I12145,g158,I12143);
  ND2 NAND2_241(g7596,I12127,I12128);
  ND2 NAND2_242(I13302,g8162,I13300);
  ND2 NAND2_243(I5502,g1007,I5500);
  ND2 NAND2_244(I9574,g5608,g818);
  ND2 NAND2_245(g3273,I6448,I6449);
  ND2 NAND2_246(I8670,g4831,I8669);
  ND2 NAND2_247(I7035,g1868,I7033);
  ND2 NAND2_248(I15453,g10051,I15451);
  ND2 NAND2_249(I8625,g4267,I8624);
  ND2 NAND2_250(I7876,g4109,I7875);
  ND2 NAND2_251(I14203,g8825,I14202);
  ND2 NAND2_252(I15607,g10149,g10144);
  ND2 NAND2_253(g2274,I5324,I5325);
  ND2 NAND2_254(I8740,g1121,I8738);
  ND2 NAND2_255(I17296,g11373,I17295);
  ND2 NAND2_256(g10507,g10434,g5859);
  ND2 NAND2_257(g2325,g611,g617);
  ND2 NAND2_258(I8606,g506,I8604);
  ND2 NAND2_259(I12087,g1470,I12085);
  ND2 NAND2_260(I13249,g1891,I13248);
  ND2 NAND2_261(I13248,g1891,g8148);
  ND2 NAND2_262(I13552,g668,g8262);
  ND2 NAND2_263(g2106,I4979,I4980);
  ND2 NAND2_264(I12069,g139,I12067);
  ND2 NAND2_265(g9204,g6019,g8942);
  ND2 NAND2_266(I12068,g7116,I12067);
  ND2 NAND2_267(I17503,g11475,g7603);
  ND2 NAND2_268(I7877,g810,I7875);
  ND2 NAND2_269(I5165,g1508,I5164);
  ND2 NAND2_270(g6740,g6131,g2550);
  ND2 NAND2_271(I6289,g981,I6287);
  ND2 NAND2_272(I6777,g2892,g650);
  ND2 NAND2_273(g5171,I8562,I8563);
  ND2 NAND2_274(I15891,g853,I15890);
  ND2 NAND2_275(I13090,g8006,I13089);
  ND2 NAND2_276(g11474,I17460,I17461);
  ND4 NAND4_7(g7942,g7395,g6847,g7380,g7369);
  ND2 NAND2_277(I5538,g1270,g1023);
  ND2 NAND2_278(I7563,g3533,I7562);
  ND2 NAND2_279(I13513,g686,g8248);
  ND2 NAND2_280(g2107,I4986,I4987);
  ND2 NAND2_281(g2223,I5203,I5204);
  ND2 NAND2_282(I13505,g677,I13504);
  ND2 NAND2_283(I6209,g802,I6207);
  ND2 NAND2_284(I12086,g6980,I12085);
  ND2 NAND2_285(I8545,g486,I8543);
  ND2 NAND2_286(I8180,g1786,I8178);
  ND2 NAND2_287(g2115,I5014,I5015);
  ND2 NAND2_288(I8591,g501,I8589);
  ND2 NAND2_289(I10931,g6395,I10930);
  ND2 NAND2_290(I17402,g11416,I17400);
  ND2 NAND2_291(g8307,I13294,I13295);
  ND2 NAND2_292(I12144,g7089,I12143);
  ND2 NAND2_293(I10520,g6231,I10519);
  ND2 NAND2_294(I5263,g456,g461);
  ND2 NAND2_295(g8757,g8599,g4401);
  ND2 NAND2_296(I6714,g2961,g201);
  ND2 NAND2_297(I14211,g599,I14209);
  ND2 NAND2_298(I8515,g3513,I8513);
  ND2 NAND2_299(g2272,I5316,I5317);
  ND2 NAND2_300(I9946,g5233,g1796);
  ND2 NAND2_301(I8750,g4613,g1125);
  ND2 NAND2_302(I5605,g1149,I5604);
  ND2 NAND2_303(g8880,I14203,I14204);
  ND2 NAND2_304(I16051,g837,g10371);
  ND2 NAND2_305(I16072,g845,g10373);
  ND2 NAND2_306(g10440,g10360,g6037);
  ND2 NAND2_307(g8612,I13858,I13859);
  ND2 NAND2_308(I15872,g2713,I15870);
  ND2 NAND2_309(I8528,g4879,I8527);
  ND2 NAND2_310(g8629,I13901,I13902);
  ND4 NAND4_8(g8542,g2571,g1828,g1814,g8390);
  ND2 NAND2_311(I9947,g5233,I9946);
  ND2 NAND2_312(I6838,g806,I6836);
  ND2 NAND2_313(g7583,I12068,I12069);
  ND2 NAND2_314(g4803,g3664,g2356);
  ND2 NAND2_315(I17307,g11377,I17305);
  ND2 NAND2_316(g4538,g3475,g2399);
  ND2 NAND2_317(I15452,g10058,I15451);
  ND2 NAND2_318(I13857,g8538,g1448);
  ND2 NAND2_319(I14202,g8825,g591);
  ND2 NAND2_320(I13765,g731,g8417);
  ND2 NAND2_321(g2260,I5296,I5297);
  ND4 NAND4_9(g7986,g7011,g6995,g6984,g7550);
  ND2 NAND2_322(g5226,I8670,I8671);
  ND2 NAND2_323(g8512,g3723,g8366);
  ND2 NAND2_324(I16046,g10370,I16044);
  ND2 NAND2_325(I13504,g677,g8247);
  ND2 NAND2_326(g10447,g10363,g5360);
  ND2 NAND2_327(g2167,I5105,I5106);
  ND2 NAND2_328(I8804,g4677,I8803);
  ND2 NAND2_329(g10472,I16016,I16017);
  ND2 NAND2_330(I17487,g11474,I17485);
  ND2 NAND2_331(I4995,g416,g309);
  ND2 NAND2_332(I12093,g6944,I12092);
  ND4 NAND4_10(g7987,g7011,g6995,g7562,g6974);
  ND2 NAND2_333(g5227,I8677,I8678);
  ND2 NAND2_334(I5126,g1386,g1389);
  ND2 NAND2_335(g2321,I5372,I5373);
  ND2 NAND2_336(g7547,I11974,I11975);
  ND2 NAND2_337(I17306,g11381,I17305);
  ND3 NAND3_4(g6548,g6132,g6124,g6122);
  ND2 NAND2_338(I11995,g7107,g127);
  ND2 NAND2_339(I7225,g1781,I7223);
  ND2 NAND2_340(I11261,g6775,g826);
  ND3 NAND3_5(g8843,g8542,g8757,g8545);
  ND2 NAND2_341(g2938,I6110,I6111);
  ND2 NAND2_342(I4942,g396,I4941);
  ND2 NAND2_343(g10394,I15899,I15900);
  ND2 NAND2_344(g8549,g5527,g8390);
  ND2 NAND2_345(g3070,g2016,g1206);
  ND2 NAND2_346(I4954,g401,g327);
  ND2 NAND2_347(I5023,g995,g1275);
  ND2 NAND2_348(g10446,g10443,g5350);
  ND2 NAND2_349(I16081,g10374,I16079);
  ND2 NAND2_350(I8641,g4278,I8640);
  ND2 NAND2_351(I6178,g197,I6176);
  ND2 NAND2_352(I12075,g7098,I12074);
  ND2 NAND2_353(I5127,g1386,I5126);
  ND2 NAND2_354(I5451,g991,I5449);
  ND2 NAND2_355(g4168,I7322,I7323);
  ND2 NAND2_356(I6288,g2091,I6287);
  ND2 NAND2_357(I8179,g3685,I8178);
  ND2 NAND2_358(I4912,g318,I4910);
  ND2 NAND2_359(I6805,g3268,g471);
  ND3 NAND3_6(g3766,g2439,g3222,g2493);
  ND2 NAND2_360(g3087,I6288,I6289);
  ND2 NAND2_361(I17486,g11384,I17485);
  ND2 NAND2_362(I4929,g391,I4928);
  ND2 NAND2_363(I15890,g853,g10286);
  ND2 NAND2_364(I16331,g10616,I16330);
  ND2 NAND2_365(I9575,g5608,I9574);
  ND2 NAND2_366(I13887,g8532,I13886);
  ND2 NAND2_367(g5308,I8787,I8788);
  ND2 NAND2_368(I13529,g704,g8253);
  ND2 NAND2_369(I6208,g2534,I6207);
  ND2 NAND2_370(g5217,I8641,I8642);
  ND2 NAND2_371(I5316,g1032,I5315);
  ND2 NAND2_372(g2111,I5006,I5007);
  ND2 NAND2_373(g10366,g10285,g5392);
  ND2 NAND2_374(I5034,g1015,g1019);
  ND2 NAND2_375(I13869,g1403,I13867);
  ND2 NAND2_376(I13868,g8523,I13867);
  ND2 NAND2_377(I15999,g10423,g2683);
  ND2 NAND2_378(I13259,g1900,I13258);
  ND4 NAND4_11(g3261,g2229,g2222,g2211,g2202);
  ND2 NAND2_379(g10481,I16073,I16074);
  ND2 NAND2_380(g2180,I5136,I5137);
  ND3 NAND3_7(g4976,g2310,g4604,g3807);
  ND2 NAND2_381(g8506,g3475,g8366);
  ND2 NAND2_382(g2380,I5460,I5461);
  ND2 NAND2_383(I13258,g1900,g8153);
  ND2 NAND2_384(I5013,g1007,g1011);
  ND2 NAND2_385(g5196,I8605,I8606);
  ND2 NAND2_386(I10930,g6395,g5555);
  ND2 NAND2_387(I6770,g3257,g382);
  ND2 NAND2_388(g11449,I17401,I17402);
  ND2 NAND2_389(g11448,I17394,I17395);
  ND2 NAND2_390(I15717,g10231,I15716);
  ND2 NAND2_391(I5317,g1027,I5315);
  ND2 NAND2_392(I14210,g8824,I14209);
  ND2 NAND2_393(I17569,g1610,I17567);
  ND2 NAND2_394(I13878,g1444,I13876);
  ND2 NAND2_395(g8545,g3710,g8390);
  ND2 NAND2_396(g2515,I5605,I5606);
  ND2 NAND2_397(I14443,g8970,I14442);
  ND2 NAND2_398(g7557,I11996,I11997);
  ND2 NAND2_399(g8180,I13090,I13091);
  ND2 NAND2_400(I14279,g1828,I14277);
  ND2 NAND2_401(I17568,g11496,I17567);
  ND2 NAND2_402(I13886,g8532,g1440);
  ND2 NAND2_403(I7322,g3047,I7321);
  ND2 NAND2_404(I6990,g986,I6988);
  ND2 NAND2_405(I14278,g8847,I14277);
  ND2 NAND2_406(I7033,g3089,g1868);
  ND2 NAND2_407(I9006,g4492,g1791);
  ND2 NAND2_408(g8507,g3738,g8366);
  ND2 NAND2_409(I5460,g1240,I5459);
  ND2 NAND2_410(g4588,g3440,g2745);
  ND2 NAND2_411(I4986,g999,I4985);
  ND3 NAND3_8(g3247,g1828,g2564,g2571);
  ND2 NAND2_412(I8651,g4824,I8650);
  ND2 NAND2_413(I13545,g713,I13544);
  ND2 NAND2_414(g8628,I13894,I13895);
  ND2 NAND2_415(I6138,g378,I6136);
  ND2 NAND2_416(I12074,g7098,g174);
  ND2 NAND2_417(g8630,I13908,I13909);
  ND2 NAND2_418(I13078,g7963,I13076);
  ND2 NAND2_419(I6109,g2205,g1494);
  ND2 NAND2_420(g8300,I13259,I13260);
  ND2 NAND2_421(I5501,g1255,I5500);
  ND2 NAND2_422(I17586,g11515,I17584);
  ND2 NAND2_423(I12092,g6944,g1490);
  ND2 NAND2_424(I13901,g8520,I13900);
  ND2 NAND2_425(I8795,g4672,g1145);
  ND2 NAND2_426(I6201,g766,I6199);
  ND2 NAND2_427(I14217,g8826,I14216);
  ND2 NAND2_428(I9007,g4492,I9006);
  ND2 NAND2_429(I13561,g8263,I13559);
  ND2 NAND2_430(I15716,g10231,g10229);
  ND2 NAND2_431(I6449,g1776,I6447);
  ND2 NAND2_432(I13295,g8161,I13293);
  ND2 NAND2_433(I4987,g1003,I4985);
  ND2 NAND2_434(I6715,g2961,I6714);
  ND2 NAND2_435(I17493,g11475,I17492);
  ND2 NAND2_436(I12215,g7061,I12214);
  ND2 NAND2_437(g2372,I5450,I5451);
  ND2 NAND2_438(g7062,I11262,I11263);
  ND2 NAND2_439(g2988,I6225,I6226);
  ND2 NAND2_440(I13309,g617,I13307);
  ND2 NAND2_441(g8839,g8750,g4401);
  ND2 NAND2_442(g2555,I5676,I5677);
  ND2 NAND2_443(g3662,I6826,I6827);
  ND2 NAND2_444(I13308,g8190,I13307);
  ND2 NAND2_445(g2792,I5879,I5880);
  ND2 NAND2_446(g4117,g3041,g3061);
  ND2 NAND2_447(I8543,g4218,g486);
  ND2 NAND2_448(g11549,I17585,I17586);
  ND2 NAND2_449(I6881,g1351,I6879);
  ND2 NAND2_450(I12138,g131,I12136);
  ND2 NAND2_451(I8729,g4605,I8728);
  ND2 NAND2_452(I14216,g8826,g605);
  ND2 NAND2_453(g10384,I15871,I15872);
  ND2 NAND2_454(I13260,g8153,I13258);
  ND2 NAND2_455(g2776,I5866,I5867);
  ND2 NAND2_456(I8513,g4873,g3513);
  ND2 NAND2_457(I13559,g722,g8263);
  ND2 NAND2_458(I8178,g3685,g1786);
  ND2 NAND2_459(g3631,I6793,I6794);
  ND2 NAND2_460(I6487,g2306,g1227);
  ND2 NAND2_461(I16080,g849,I16079);
  ND2 NAND2_462(I13893,g8529,g1436);
  ND2 NAND2_463(I12115,g162,I12113);
  ND2 NAND2_464(I6748,g1453,I6746);
  ND2 NAND2_465(I13544,g713,g8259);
  ND2 NAND2_466(I5484,g1250,g1011);
  ND2 NAND2_467(I4928,g391,g321);
  ND2 NAND2_468(I6226,g1346,I6224);
  ND2 NAND2_469(I8805,g1113,I8803);
  ND2 NAND2_470(I4930,g321,I4928);
  ND2 NAND2_471(I15880,g2719,I15878);
  ND2 NAND2_472(I14265,g1814,I14263);
  ND2 NAND2_473(I16031,g829,I16030);
  ND2 NAND2_474(g3585,I6747,I6748);
  ND4 NAND4_12(g3041,g2364,g2399,g2374,g2382);
  ND2 NAND2_475(g8933,I14271,I14272);
  ND2 NAND2_476(I16330,g10616,g4997);
  ND2 NAND2_477(I13267,g8154,I13265);
  ND2 NAND2_478(I13294,g1882,I13293);
  ND2 NAND2_479(g10231,I15616,I15617);
  ND2 NAND2_480(I14442,g8970,g1834);
  ND2 NAND2_481(I6793,g2959,I6792);
  ND2 NAND2_482(I4966,g330,I4964);
  ND2 NAND2_483(I8752,g1125,I8750);
  ND2 NAND2_484(I15432,g10044,I15430);
  ND2 NAND2_485(I12214,g7061,g2518);
  ND2 NAND2_486(g10511,g10438,g6032);
  ND2 NAND2_487(g3011,g591,g2382);
  ND2 NAND2_488(g5103,I8480,I8481);
  ND2 NAND2_489(I16087,g861,I16086);
  ND2 NAND2_490(g3734,g3039,g599);
  ND2 NAND2_491(I6664,g2792,g2776);
  ND2 NAND2_492(g8882,I14217,I14218);
  ND2 NAND2_493(I4955,g401,I4954);
  ND2 NAND2_494(I8786,g4639,g1141);
  ND3 NAND3_9(g3992,g2571,g2550,g2990);
  ND2 NAND2_495(g10480,I16066,I16067);
  ND2 NAND2_496(I11915,g6935,I11914);
  ND2 NAND2_497(I8770,g4619,g1133);
  ND2 NAND2_498(I5516,g1260,g1019);
  ND2 NAND2_499(g8541,g4001,g8390);
  ND2 NAND2_500(I6188,g466,I6186);
  ND2 NAND2_501(g5147,I8544,I8545);
  ND3 NAND3_10(g8744,g8617,g6509,g6971);
  ND2 NAND2_502(I5892,g750,I5891);
  ND2 NAND2_503(g8558,I13766,I13767);
  ND2 NAND2_504(I15258,g9980,I15256);
  ND2 NAND2_505(I13266,g1909,I13265);
  ND2 NAND2_506(I8787,g4639,I8786);
  ND2 NAND2_507(I6826,g3281,I6825);
  ND2 NAND2_508(I17283,g11357,I17281);
  ND3 NAND3_11(g5013,g4749,g3247,g3205);
  ND2 NAND2_509(I17492,g11475,g3623);
  ND2 NAND2_510(g8511,g5277,g8366);
  ND2 NAND2_511(I16079,g849,g10374);
  ND2 NAND2_512(I5035,g1015,I5034);
  ND2 NAND2_513(I5517,g1260,I5516);
  ND2 NAND2_514(I7223,g2981,g1781);
  ND2 NAND2_515(I16086,g861,g10375);
  ND2 NAND2_516(g5317,I8796,I8797);
  ND2 NAND2_517(I15879,g10359,I15878);
  ND2 NAND2_518(I15878,g10359,g2719);
  ND2 NAND2_519(I12114,g7093,I12113);
  ND2 NAND2_520(I12107,g7113,I12106);
  ND2 NAND2_521(g2500,g178,g182);
  ND2 NAND2_522(I15994,g2677,I15992);
  ND4 NAND4_13(g7934,g7395,g6847,g7279,g7369);
  ND2 NAND2_523(g10469,g10430,g5999);
  ND2 NAND2_524(I14264,g8843,I14263);
  ND2 NAND2_525(I6448,g2264,I6447);
  ND2 NAND2_526(I13285,g8159,I13283);
  ND2 NAND2_527(g10468,I16000,I16001);
  ND2 NAND2_528(I6827,g770,I6825);
  ND2 NAND2_529(g8623,I13877,I13878);
  ND2 NAND2_530(I13900,g8520,g1428);
  ND2 NAND2_531(g2795,I5892,I5893);
  ND2 NAND2_532(I8575,g4234,g496);
  ND2 NAND2_533(I14209,g8824,g599);
  ND2 NAND2_534(I13560,g722,I13559);
  ND2 NAND2_535(I8715,g4601,g4052);
  ND2 NAND2_536(I8604,g4259,g506);
  ND2 NAND2_537(I16017,g2695,I16015);
  ND2 NAND2_538(I4941,g396,g324);
  ND2 NAND2_539(g2205,I5165,I5166);
  ND3 NAND3_12(g3753,g2382,g2364,g2800);
  ND2 NAND2_540(I6467,g23,g2479);
  ND2 NAND2_541(I14614,g611,I14612);
  ND2 NAND2_542(g2104,I4965,I4966);
  ND2 NAND2_543(g2099,I4942,I4943);
  ND2 NAND2_544(I16023,g10426,g2701);
  ND2 NAND2_545(g10479,I16059,I16060);
  ND3 NAND3_13(g8737,g2317,g4921,g8688);
  ND2 NAND2_546(g5942,I9575,I9576);
  ND2 NAND2_547(g10478,I16052,I16053);
  ND2 NAND2_548(I12004,g153,I12002);
  ND2 NAND2_549(I4911,g386,I4910);
  ND2 NAND2_550(I11914,g6935,g1494);
  ND2 NAND2_551(g7960,g7409,g5573);
  ND2 NAND2_552(I5295,g794,g798);
  ND2 NAND2_553(I12106,g7113,g135);
  ND2 NAND2_554(I8728,g4605,g1117);
  ND2 NAND2_555(g3681,I6837,I6838);
  ND2 NAND2_556(I11907,g6967,g1474);
  ND2 NAND2_557(I13907,g8526,g1432);
  ND2 NAND2_558(I8730,g1117,I8728);
  ND2 NAND2_559(g8551,g3967,g8390);
  ND2 NAND2_560(I4980,g333,I4978);
  ND2 NAND2_561(g2961,I6177,I6178);
  ND2 NAND2_562(g6019,g617,g4921);
  ND2 NAND2_563(I16016,g10425,I16015);
  ND2 NAND2_564(I11935,g7004,g1458);
  ND2 NAND2_565(I8678,g1027,I8676);
  ND2 NAND2_566(I17051,g10923,g11249);
  ND2 NAND2_567(g4482,I7864,I7865);
  ND2 NAND2_568(g7592,I12107,I12108);
  ND2 NAND2_569(g3460,I6665,I6666);
  ND4 NAND4_14(g7932,g7395,g6847,g7279,g7273);
  ND2 NAND2_570(g7624,I12215,I12216);
  ND4 NAND4_15(g7953,g7395,g7390,g7380,g7369);
  ND2 NAND2_571(g8414,I13553,I13554);
  ND2 NAND2_572(I6168,g153,I6166);
  ND2 NAND2_573(I5229,g182,g148);
  ND2 NAND2_574(I6772,g382,I6770);
  ND2 NAND2_575(I16030,g829,g10368);
  ND2 NAND2_576(I13284,g1927,I13283);
  ND2 NAND2_577(I16065,g10428,g2765);
  ND2 NAND2_578(g2947,I6137,I6138);
  ND2 NAND2_579(I7321,g3047,g1231);
  ND2 NAND2_580(g2437,I5529,I5530);
  ND2 NAND2_581(g2102,I4955,I4956);
  ND2 NAND2_582(I17282,g11360,I17281);
  ND2 NAND2_583(I5620,g1771,I5618);
  ND2 NAND2_584(I8664,g476,I8662);
  ND2 NAND2_585(g7524,I11915,I11916);
  ND2 NAND2_586(g7717,g6863,g3206);
  ND2 NAND2_587(I16467,g10716,g10518);
  ND2 NAND2_588(I4972,g991,I4971);
  ND2 NAND2_589(I13554,g8262,I13552);
  ND2 NAND2_590(I16037,g10427,g2707);
  ND2 NAND2_591(g8302,I13273,I13274);
  ND2 NAND2_592(I4943,g324,I4941);
  ND2 NAND2_593(I5485,g1250,I5484);
  ND2 NAND2_594(g5527,g3978,g4749);
  ND2 NAND2_595(I10509,g786,I10507);
  ND2 NAND2_596(g7599,I12144,I12145);
  ND2 NAND2_597(I10508,g6221,I10507);
  ND2 NAND2_598(I6126,g1419,I6124);
  ND2 NAND2_599(I8671,g814,I8669);
  ND2 NAND2_600(I6760,g2943,g1448);
  ND2 NAND2_601(g3626,I6778,I6779);
  ND2 NAND2_602(I11973,g7001,g1462);
  ND2 NAND2_603(g2389,I5469,I5470);
  ND2 NAND2_604(I15617,g10153,I15615);
  ND2 NAND2_605(g5277,g3734,g4538);
  ND2 NAND2_606(I5005,g421,g312);
  ND2 NAND2_607(I6779,g650,I6777);
  ND2 NAND2_608(I6665,g2792,I6664);
  ND2 NAND2_609(I8589,g4251,g501);
  ND2 NAND2_610(g8412,I13545,I13546);
  ND2 NAND2_611(g2963,I6187,I6188);
  ND2 NAND2_612(I12045,g6951,g1486);
  ND2 NAND2_613(I16053,g10371,I16051);
  ND2 NAND2_614(g2109,I4996,I4997);
  ND2 NAND2_615(g11418,I17306,I17307);
  ND2 NAND2_616(I13539,g8157,I13537);
  ND2 NAND2_617(g10475,I16031,I16032);
  ND2 NAND2_618(I5324,g1336,I5323);
  ND2 NAND2_619(I13538,g658,I13537);
  ND2 NAND2_620(I5469,g1245,I5468);
  ND2 NAND2_621(I5540,g1023,I5538);
  ND2 NAND2_622(I17505,g7603,I17503);
  ND2 NAND2_623(I11241,g6760,g790);
  ND2 NAND2_624(I8803,g4677,g1113);
  ND2 NAND2_625(I12061,g6961,I12060);
  ND2 NAND2_626(I8780,g1137,I8778);
  ND3 NAND3_14(g8745,g8617,g6517,g6964);
  ND2 NAND2_627(I4979,g411,I4978);
  ND2 NAND2_628(g8109,g5052,g7853);
  ND2 NAND2_629(g8309,I13308,I13309);
  ND2 NAND2_630(g6758,I10770,I10771);
  ND2 NAND2_631(I16009,g2689,I16007);
  ND2 NAND2_632(I15616,g10043,I15615);
  ND2 NAND2_633(I8662,g4286,g476);
  ND2 NAND2_634(I16008,g10424,I16007);
  ND2 NAND2_635(I13515,g8248,I13513);
  ND2 NAND2_636(I13991,g622,I13990);
  ND2 NAND2_637(g11276,I17052,I17053);
  ND2 NAND2_638(I15900,g10287,I15898);
  ND2 NAND2_639(g2419,I5501,I5502);
  ND2 NAND2_640(I16074,g10373,I16072);
  ND2 NAND2_641(I10769,g5944,g1801);
  ND2 NAND2_642(I7323,g1231,I7321);
  ND2 NAND2_643(g7978,g7697,g3038);
  ND2 NAND2_644(I7875,g4109,g810);
  ND2 NAND2_645(I8562,g4227,I8561);
  ND2 NAND2_646(I15892,g10286,I15890);
  ND2 NAND2_647(g3771,I6989,I6990);
  ND2 NAND2_648(I8605,g4259,I8604);
  ND2 NAND2_649(g10153,I15452,I15453);
  ND2 NAND2_650(g5295,I8762,I8763);
  ND2 NAND2_651(I8751,g4613,I8750);
  ND2 NAND2_652(I15907,g6899,I15906);
  ND2 NAND2_653(I5136,g521,I5135);
  ND2 NAND2_654(I11263,g826,I11261);
  ND2 NAND2_655(I14204,g591,I14202);
  ND2 NAND2_656(g8881,I14210,I14211);
  ND2 NAND2_657(g2105,I4972,I4973);
  ND3 NAND3_15(g5557,g4538,g3071,g3011);
  ND2 NAND2_658(I5230,g182,I5229);
  ND2 NAND2_659(I8669,g4831,g814);
  ND2 NAND2_660(g10474,I16024,I16025);
  ND2 NAND2_661(I8772,g1133,I8770);
  ND2 NAND2_662(g2445,I5539,I5540);
  ND2 NAND2_663(g8006,g5552,g7717);
  ND2 NAND2_664(I10932,g5555,I10930);
  ND2 NAND2_665(I17504,g11475,I17503);
  ND2 NAND2_666(I5137,g525,I5135);
  ND2 NAND2_667(g8305,I13284,I13285);
  ND2 NAND2_668(I5891,g750,g2057);
  ND2 NAND2_669(I13273,g1918,I13272);
  ND2 NAND2_670(I8480,g4455,I8479);
  ND2 NAND2_671(g4144,g2160,g3044);
  ND2 NAND2_672(I15906,g6899,g10302);
  ND2 NAND2_673(I5342,g315,I5341);
  ND2 NAND2_674(I13514,g686,I13513);
  ND2 NAND2_675(g8407,I13522,I13523);
  ND2 NAND2_676(g4088,I7224,I7225);
  ND2 NAND2_677(g4488,I7876,I7877);
  ND2 NAND2_678(g7598,I12137,I12138);
  ND3 NAND3_16(g3222,g2557,g1814,g1834);
  ND2 NAND2_679(I16052,g837,I16051);
  ND2 NAND2_680(I12127,g7103,I12126);
  ND2 NAND2_681(g10483,I16087,I16088);
  ND2 NAND2_682(g8415,I13560,I13561);
  ND2 NAND2_683(g11415,I17289,I17290);
  ND2 NAND2_684(g6573,I10508,I10509);
  ND2 NAND2_685(I5676,g1218,I5675);
  ND2 NAND2_686(I6778,g2892,I6777);
  ND2 NAND2_687(g9413,I14613,I14614);
  ND2 NAND2_688(I8779,g4630,I8778);
  ND2 NAND2_689(I5592,g1696,I5591);
  ND4 NAND4_16(g8502,g2382,g605,g591,g8366);
  ND2 NAND2_690(I15609,g10144,I15607);
  ND2 NAND2_691(I15608,g10149,I15607);
  ND3 NAND3_17(g3071,g605,g2374,g2382);
  ND2 NAND2_692(g10509,g10436,g6023);
  ND2 NAND2_693(I17461,g11448,I17459);
  ND2 NAND2_694(I13506,g8247,I13504);
  ND2 NAND2_695(I5468,g1245,g999);
  ND2 NAND2_696(g5219,I8651,I8652);
  ND2 NAND2_697(I5677,g1223,I5675);
  ND3 NAND3_18(g8826,g8739,g8737,g8648);
  ND2 NAND2_698(I17393,g11415,g11414);
  ND2 NAND2_699(I5866,g2107,I5865);
  ND2 NAND2_700(I12126,g7103,g170);
  ND2 NAND2_701(I4978,g411,g333);
  ND2 NAND2_702(g7587,I12086,I12087);
  ND2 NAND2_703(g5286,I8751,I8752);
  ND2 NAND2_704(g8308,I13301,I13302);
  ND2 NAND2_705(I7864,g4099,I7863);
  ND2 NAND2_706(I11981,g6957,I11980);
  ND2 NAND2_707(I12060,g6961,g1478);
  ND2 NAND2_708(g5225,I8663,I8664);
  ND2 NAND2_709(g11538,I17568,I17569);
  ND2 NAND2_710(I13767,g8417,I13765);
  ND2 NAND2_711(g10396,I15907,I15908);
  ND2 NAND2_712(I11262,g6775,I11261);
  ND2 NAND2_713(I13990,g622,g8688);
  ND2 NAND2_714(I6224,g2544,g1346);
  ND2 NAND2_715(I5867,g2105,I5865);
  ND2 NAND2_716(g2493,g1834,g1840);
  ND2 NAND2_717(I5893,g2057,I5891);
  ND3 NAND3_19(g3062,g2369,g591,g611);
  ND2 NAND2_718(I13521,g695,g8249);
  ND2 NAND2_719(I5186,g1515,I5184);
  ND2 NAND2_720(I6771,g3257,I6770);
  ND2 NAND2_721(I5325,g1341,I5323);
  ND2 NAND2_722(I17459,g11449,g11448);
  ND2 NAND2_723(I9557,g5598,g782);
  ND2 NAND2_724(g11414,I17282,I17283);
  ND2 NAND2_725(I12067,g7116,g139);
  ND2 NAND2_726(I12094,g1490,I12092);
  ND2 NAND2_727(I4964,g406,g330);
  ND2 NAND2_728(I13272,g1918,g8158);
  ND2 NAND2_729(I9948,g1796,I9946);
  ND2 NAND2_730(g10302,I15717,I15718);
  ND2 NAND2_731(I16332,g4997,I16330);
  ND2 NAND2_732(I5106,g435,I5104);
  ND2 NAND2_733(g8847,g8760,g8683);
  ND2 NAND2_734(g2257,I5283,I5284);
  ND2 NAND2_735(I12019,g7119,g166);
  ND2 NAND2_736(I15441,g10035,g10122);
  ND2 NAND2_737(I11997,g127,I11995);
  ND2 NAND2_738(I8739,g4607,I8738);
  ND2 NAND2_739(I5461,g1003,I5459);
  ND2 NAND2_740(I13766,g731,I13765);
  ND2 NAND2_741(I8479,g4455,g3530);
  ND2 NAND2_742(I17295,g11373,g11369);
  ND2 NAND2_743(I14271,g8840,I14270);
  ND2 NAND2_744(I4971,g991,g995);
  ND2 NAND2_745(g8301,I13266,I13267);
  ND2 NAND2_746(I6110,g2205,I6109);
  ND2 NAND2_747(g10482,I16080,I16081);
  ND2 NAND2_748(g10779,I16468,I16469);
  ND2 NAND2_749(I6762,g1448,I6760);
  ND2 NAND2_750(I17289,g11366,I17288);
  ND2 NAND2_751(I5315,g1032,g1027);
  ND2 NAND2_752(I17288,g11366,g11363);
  ND2 NAND2_753(I13859,g1448,I13857);
  ND2 NAND2_754(g7548,I11981,I11982);
  ND2 NAND2_755(I13858,g8538,I13857);
  ND2 NAND2_756(I11996,g7107,I11995);
  ND3 NAND3_20(g8743,g8617,g6971,g6964);
  ND2 NAND2_757(I5880,g2115,I5878);
  ND2 NAND2_758(g10513,g10441,g5345);
  ND2 NAND2_759(g8411,I13538,I13539);
  ND2 NAND2_760(I8626,g511,I8624);
  ND2 NAND2_761(g10505,g10432,g5938);
  ND2 NAND2_762(I5612,g1280,I5611);
  ND2 NAND2_763(g4821,I8179,I8180);
  ND2 NAND2_764(I12076,g174,I12074);
  ND2 NAND2_765(I12085,g6980,g1470);
  ND2 NAND2_766(g7567,I12020,I12021);
  ND2 NAND2_767(I5128,g1389,I5126);
  ND2 NAND2_768(I6489,g1227,I6487);
  ND2 NAND2_769(g7593,I12114,I12115);
  ND2 NAND2_770(I8778,g4630,g1137);
  ND2 NAND2_771(g10149,I15442,I15443);
  ND2 NAND2_772(I13902,g1428,I13900);
  ND2 NAND2_773(I13301,g1936,I13300);
  ND2 NAND2_774(g3215,g2564,g1822);
  ND4 NAND4_17(g7996,g7011,g7574,g7562,g6974);
  ND2 NAND2_775(I4985,g999,g1003);
  ND2 NAND2_776(I14444,g1834,I14442);
  ND4 NAND4_18(g8000,g7011,g7574,g7562,g7550);
  ND2 NAND2_777(I5166,g1499,I5164);
  ND2 NAND2_778(I17460,g11449,I17459);
  ND2 NAND2_779(g3008,g2444,g878);
  ND2 NAND2_780(I6836,g3287,g806);
  ND2 NAND2_781(I5529,g1265,I5528);
  ND2 NAND2_782(g10229,I15608,I15609);
  ND2 NAND2_783(I13661,g8322,I13659);
  ND2 NAND2_784(I13895,g1436,I13893);
  ND2 NAND2_785(g2303,I5342,I5343);
  ND2 NAND2_786(I12039,g6990,I12038);
  ND2 NAND2_787(g5592,I9007,I9008);
  ND2 NAND2_788(I12038,g6990,g1466);
  ND2 NAND2_789(g3322,I6488,I6489);
  ND2 NAND2_790(I8561,g4227,g491);
  ND2 NAND2_791(I8527,g4879,g481);
  ND2 NAND2_792(I12143,g7089,g158);
  ND2 NAND2_793(I5619,g1766,I5618);
  ND2 NAND2_794(g10386,I15879,I15880);
  ND2 NAND2_795(I11980,g6957,g1482);
  ND2 NAND2_796(I6837,g3287,I6836);
  ND2 NAND2_797(I4973,g995,I4971);
  ND2 NAND2_798(I13888,g1440,I13886);
  ND2 NAND2_799(g7558,I12003,I12004);
  ND2 NAND2_800(I17494,g3623,I17492);
  ND2 NAND2_801(g11491,I17493,I17494);
  ND2 NAND2_802(I16045,g833,I16044);
  ND2 NAND2_803(I7684,g1023,I7683);
  ND2 NAND2_804(g4130,g3044,g2518);
  ND2 NAND2_805(I8771,g4619,I8770);
  ND2 NAND2_806(I13546,g8259,I13544);
  ND2 NAND2_807(I13089,g8006,g1840);
  ND2 NAND2_808(g2117,I5024,I5025);
  ND2 NAND2_809(g5119,I8514,I8515);
  ND2 NAND2_810(g5319,I8804,I8805);
  ND2 NAND2_811(I15899,g857,I15898);
  ND2 NAND2_812(I5606,g1153,I5604);
  ND2 NAND2_813(I15898,g857,g10287);
  ND2 NAND2_814(I16032,g10368,I16030);
  ND2 NAND2_815(I17401,g11418,I17400);
  ND2 NAND2_816(I13659,g1945,g8322);
  ND2 NAND2_817(I8738,g4607,g1121);
  ND2 NAND2_818(I13250,g8148,I13248);
  ND2 NAND2_819(I15718,g10229,I15716);
  ND2 NAND2_820(I9008,g1791,I9006);
  ND2 NAND2_821(I6176,g2177,g197);
  ND2 NAND2_822(I7865,g774,I7863);
  ND2 NAND2_823(g5274,I8729,I8730);
  ND2 NAND2_824(I5341,g315,g426);
  ND2 NAND2_825(I17305,g11381,g11377);
  ND2 NAND2_826(I17053,g11249,I17051);
  ND2 NAND2_827(g5125,I8528,I8529);
  ND2 NAND2_828(I12216,g2518,I12214);
  ND2 NAND2_829(I6225,g2544,I6224);
  ND2 NAND2_830(I5879,g2120,I5878);
  ND2 NAND2_831(g3221,g1834,g2564);
  ND2 NAND2_832(I14270,g8840,g1822);
  ND2 NAND2_833(I6124,g2215,g1419);
  ND2 NAND2_834(I6324,g1864,I6322);
  ND2 NAND2_835(I13867,g8523,g1403);
  ND2 NAND2_836(I13894,g8529,I13893);
  ND2 NAND2_837(I6469,g2479,I6467);
  ND2 NAND2_838(I8663,g4286,I8662);
  ND2 NAND2_839(g7523,I11908,I11909);
  ND2 NAND2_840(I6177,g2177,I6176);
  ND2 NAND2_841(g5187,I8590,I8591);
  ND2 NAND2_842(I6287,g2091,g981);
  ND2 NAND2_843(I8762,g4616,I8761);
  ND2 NAND2_844(I15871,g10358,I15870);
  ND3 NAND3_21(g8840,g8542,g8541,g8760);
  ND2 NAND2_845(g2250,I5264,I5265);
  ND2 NAND2_846(I8590,g4251,I8589);
  ND2 NAND2_847(I6199,g2525,g766);
  ND2 NAND2_848(I14218,g605,I14216);
  ND2 NAND2_849(g8190,g6027,g7978);
  ND2 NAND2_850(I5284,g762,I5282);
  ND2 NAND2_851(I17485,g11384,g11474);
  ND2 NAND2_852(I4965,g406,I4964);
  ND2 NAND2_853(I5591,g1696,g1703);
  ND2 NAND2_854(g8501,g3760,g8366);
  ND2 NAND2_855(I15451,g10058,g10051);
  ND2 NAND2_856(g8942,g8823,g4921);
  ND2 NAND2_857(I13877,g8535,I13876);
  ND2 NAND2_858(g7269,I11509,I11510);
  ND2 NAND2_859(I4996,g416,I4995);
  ND2 NAND2_860(I6144,g1976,I6143);
  ND2 NAND2_861(I17567,g11496,g1610);
  ND2 NAND2_862(g7572,I12039,I12040);
  ND2 NAND2_863(I6207,g2534,g802);
  ND2 NAND2_864(I14277,g8847,g1828);
  ND2 NAND2_865(I16059,g841,I16058);
  ND2 NAND2_866(I16025,g2701,I16023);
  ND2 NAND2_867(I8563,g491,I8561);
  ND2 NAND2_868(g3524,g3209,g3221);
  ND2 NAND2_869(I16058,g841,g10372);
  ND2 NAND2_870(I5204,g374,I5202);
  ND2 NAND2_871(I6488,g2306,I6487);
  ND4 NAND4_19(g3818,g3056,g3071,g2310,g3003);
  ND2 NAND2_872(I16044,g833,g10370);
  ND2 NAND2_873(g3717,I6880,I6881);
  ND2 NAND2_874(I13077,g1872,I13076);
  ND2 NAND2_875(g10043,I15257,I15258);
  ND2 NAND2_876(I11280,g6485,I11278);
  ND2 NAND2_877(I6825,g3281,g770);
  ND2 NAND2_878(I4997,g309,I4995);
  ND2 NAND2_879(I13300,g1936,g8162);
  ND2 NAND2_880(I5323,g1336,g1341);
  ND2 NAND2_881(I6136,g2496,g378);
  ND2 NAND2_882(g5935,I9558,I9559);
  ND2 NAND2_883(I5528,g1265,g1015);
  ND2 NAND2_884(I6806,g3268,I6805);
  ND2 NAND2_885(I5530,g1015,I5528);
  ND2 NAND2_886(g10886,g10807,g10805);
  ND2 NAND2_887(g3106,I6323,I6324);
  ND2 NAND2_888(I13876,g8535,g1444);
  ND2 NAND2_889(I6322,g2050,g1864);
  ND2 NAND2_890(g3061,g611,g2374);
  ND2 NAND2_891(g2439,g1814,g1828);
  ND4 NAND4_20(g7947,g7395,g7390,g7279,g7369);
  ND2 NAND2_892(I9576,g818,I9574);
  ND2 NAND2_893(I13660,g1945,I13659);
  ND2 NAND2_894(g3200,g1822,g2061);
  ND2 NAND2_895(g4374,I7684,I7685);
  ND2 NAND2_896(I11916,g1494,I11914);
  ND2 NAND2_897(I5372,g971,I5371);
  ND2 NAND2_898(g3003,g599,g2399);
  ND2 NAND2_899(g8627,I13887,I13888);
  ND2 NAND2_900(I5618,g1766,g1771);
  ND2 NAND2_901(I6137,g2496,I6136);
  ND2 NAND2_902(I5343,g426,I5341);
  ND2 NAND2_903(I5282,g758,g762);
  ND2 NAND2_904(I13307,g8190,g617);
  ND2 NAND2_905(I13076,g1872,g7963);
  ND2 NAND2_906(I6807,g471,I6805);
  ND2 NAND2_907(I11243,g790,I11241);
  ND2 NAND2_908(I17585,g11354,I17584);
  ND2 NAND2_909(I12137,g7110,I12136);
  ND2 NAND2_910(I7564,g654,I7562);
  ND2 NAND2_911(g2970,I6200,I6201);
  ND2 NAND2_912(g10144,I15431,I15432);
  ND2 NAND2_913(I8788,g1141,I8786);
  ND2 NAND2_914(g7054,I11242,I11243);
  ND2 NAND2_915(I17052,g10923,I17051);
  ND2 NAND2_916(g2120,I5035,I5036);
  ND2 NAND2_917(g8616,I13868,I13869);
  ND2 NAND2_918(I5202,g369,g374);
  ND2 NAND2_919(I16088,g10375,I16086);
  ND2 NAND2_920(I16024,g10426,I16023);
  ND2 NAND2_921(g11490,I17486,I17487);
  ND2 NAND2_922(I5518,g1019,I5516);
  ND3 NAND3_22(g5118,g2439,g4806,g4073);
  ND2 NAND2_923(I12021,g166,I12019);
  NR2 NOR2_0(g6392,g5859,g5938);
  NR2 NOR2_1(g5938,g2764,g4988);
  NR2 NOR2_2(g2478,g1610,g1737);
  NR2 NOR2_3(g10374,g10347,g3463);
  NR4 NOR4_0(g4278,g3800,g2593,g2586,g3776);
  NR2 NOR2_4(g10424,g10292,g4620);
  NR2 NOR2_5(g10383,g10318,g2998);
  NR2 NOR2_6(g3118,g2521,g2514);
  NR2 NOR2_7(g9815,g9392,g9367);
  NR2 NOR2_8(g11077,g10970,g10971);
  NR3 NOR3_0(g9746,g9454,g9274,g9292);
  NR3 NOR3_1(g3879,g3141,g2354,g2353);
  NR2 NOR2_9(g10285,g10276,g3566);
  NR2 NOR2_10(g11480,g11456,g4567);
  NR2 NOR2_11(g4076,g1707,g2864);
  NR2 NOR2_12(g10570,g10542,g10324);
  NR2 NOR2_13(g10239,g9317,g10179);
  NR2 NOR2_14(g10594,g10480,g10521);
  NR2 NOR2_15(g9426,g9052,g9030);
  NR2 NOR2_16(g10382,g10314,g2998);
  NR4 NOR4_1(g4672,g3501,g2669,g2662,g3479);
  NR2 NOR2_17(g5360,g2071,g4225);
  NR4 NOR4_2(g9387,g9010,g9240,g9223,I14596);
  NR2 NOR2_18(g10438,g10356,g3566);
  NR4 NOR4_3(g4613,g3077,g3491,g2662,g2655);
  NR4 NOR4_4(g9391,g9010,g9240,g9223,I14602);
  NR3 NOR3_2(g4572,g3419,g3408,g3628);
  NR3 NOR3_3(g9757,g9454,g9274,g9292);
  NR2 NOR2_19(g9416,g9052,g9030);
  NR4 NOR4_5(g9874,g9519,g9536,g9579,I15033);
  NR2 NOR2_20(g9654,g9125,g9173);
  NR4 NOR4_6(g9880,g9751,g9536,g9557,I15051);
  NR4 NOR4_7(g4873,g3292,g2593,g2586,g3776);
  NR2 NOR2_21(g2807,g22,g2320);
  NR2 NOR2_22(g10441,g10351,g3566);
  NR4 NOR4_8(g4639,g3501,g2669,g2662,g2655);
  NR2 NOR2_23(g10435,g10332,g3507);
  NR2 NOR2_24(g10849,g10739,g3903);
  NR4 NOR4_9(g9606,g9125,g9111,g9173,g9151);
  NR4 NOR4_10(g9879,g9747,g9536,g9566,I15048);
  NR2 NOR2_25(g9506,g9052,g9030);
  NR2 NOR2_26(g6155,g4974,g2864);
  NR2 NOR2_27(g6355,g6032,g6023);
  NR2 NOR2_28(g9615,g9052,g9030);
  NR2 NOR2_29(g10371,g10344,g3463);
  NR2 NOR2_30(g9591,g9125,g9151);
  NR2 NOR2_31(g10359,g10227,g4620);
  NR2 NOR2_32(g10434,g10352,g3566);
  NR2 NOR2_33(g10358,g10226,g4620);
  NR3 NOR3_4(g9750,g9454,g9274,g9292);
  NR2 NOR2_34(g10291,g10247,g3113);
  NR4 NOR4_11(g4227,g3292,g3793,g2586,g2579);
  NR4 NOR4_12(g9655,g9010,g9240,g9223,I14776);
  NR4 NOR4_13(g9410,g9010,g9240,g9223,I14607);
  NR4 NOR4_14(g9667,g9125,g9111,g9173,g9151);
  NR2 NOR2_35(g10563,g10539,g10322);
  NR2 NOR2_36(g9776,g9392,g9367);
  NR2 NOR2_37(g10324,g9317,g10244);
  NR3 NOR3_5(g4455,g3543,g3419,g3408);
  NR4 NOR4_15(g9878,g9754,g9536,g9560,I15045);
  NR2 NOR2_38(g10360,g10277,g3566);
  NR4 NOR4_16(g9882,g9742,g9536,g9563,I15057);
  NR2 NOR2_39(g10370,g10343,g3463);
  NR4 NOR4_17(g4605,g3077,g2669,g3485,g2655);
  NR2 NOR2_40(g10420,g10329,g3744);
  NR2 NOR2_41(g10562,g10483,g10529);
  NR2 NOR2_42(g10427,g10296,g4620);
  NR2 NOR2_43(g5780,g2112,g4921);
  NR2 NOR2_44(g10385,g10321,g2998);
  NR2 NOR2_45(g10376,g10323,g3113);
  NR2 NOR2_46(g10426,g10294,g4620);
  NR4 NOR4_18(g4601,g3077,g2669,g2662,g3479);
  NR2 NOR2_47(g5573,g4117,g4432);
  NR2 NOR2_48(g9808,g9392,g9367);
  NR2 NOR2_49(g5999,g2753,g4953);
  NR3 NOR3_6(g9759,g9454,g9274,g9292);
  NR2 NOR2_50(g6037,g3305,g5614);
  NR2 NOR2_51(g10287,g10275,g3463);
  NR2 NOR2_52(g5034,g3524,g4593);
  NR4 NOR4_19(g9362,g9010,g9240,g9223,I14585);
  NR4 NOR4_20(g9881,g9516,g9536,g9573,I15054);
  NR2 NOR2_53(g10443,g10353,g3566);
  NR2 NOR2_54(g10286,g10271,g3463);
  NR3 NOR3_7(g4276,g4065,g3261,g2500);
  NR4 NOR4_21(g4616,g3077,g3491,g2662,g3479);
  NR2 NOR2_55(g10363,g10355,g3566);
  NR2 NOR2_56(g2862,g2315,g2305);
  NR2 NOR2_57(g10373,g10346,g3463);
  NR2 NOR2_58(g10423,g10290,g4620);
  NR3 NOR3_8(g9758,g9454,g9274,g9292);
  NR3 NOR3_9(g9589,g9125,g9173,g9151);
  NR2 NOR2_59(g9803,g9392,g9367);
  NR2 NOR2_60(g10430,g10349,g3566);
  NR2 NOR2_61(g9421,g9052,g9030);
  NR2 NOR2_62(g10362,g10228,g3507);
  NR2 NOR2_63(g2791,g2187,g750);
  NR2 NOR2_64(g9817,g9392,g9367);
  NR4 NOR4_22(g9605,g9125,g9111,g9173,g9151);
  NR2 NOR2_65(g10372,g10345,g3463);
  NR2 NOR2_66(g9669,g9392,g9367);
  NR2 NOR2_67(g10422,g10289,g4620);
  NR2 NOR2_68(g10436,g10354,g3566);
  NR4 NOR4_23(g5556,g4787,g2695,g2299,g2031);
  NR4 NOR4_24(g4286,g3800,g2593,g3784,g2579);
  NR2 NOR2_69(g4974,g4502,g3714);
  NR2 NOR2_70(g9779,g9392,g9367);
  NR2 NOR2_71(g9423,g9052,g9030);
  NR2 NOR2_72(g5350,g4163,g4872);
  NR4 NOR4_25(g9361,g9010,g9240,g9223,I14582);
  NR4 NOR4_26(g2459,g1645,g1642,g1651,g1648);
  NR2 NOR2_73(g10381,g10310,g2998);
  NR4 NOR4_27(g4259,g3292,g3793,g3784,g3776);
  NR2 NOR2_74(g10522,g10486,g10239);
  NR2 NOR2_75(g5392,g3369,g4258);
  NR3 NOR3_10(g4122,g3291,g2410,g2538);
  NR2 NOR2_76(g6023,g2763,g4975);
  NR2 NOR2_77(g3462,g2187,g2795);
  NR4 NOR4_28(g4218,g3292,g2593,g3784,g3776);
  NR4 NOR4_29(g4267,g3800,g2593,g2586,g2579);
  NR4 NOR4_30(g4677,g3501,g2669,g3485,g2655);
  NR2 NOR2_78(g9646,g9125,g9151);
  NR2 NOR2_79(g2863,g2316,g2309);
  NR4 NOR4_31(g9616,g9010,g9240,g9223,I14751);
  NR2 NOR2_80(g6032,g3430,g5039);
  NR4 NOR4_32(g9647,g9125,g9111,g9173,g9151);
  NR2 NOR2_81(g5859,g3362,g4943);
  NR2 NOR2_82(g10433,g10330,g3507);
  NR2 NOR2_83(g10368,g10342,g3463);
  NR4 NOR4_33(g4251,g3292,g3793,g3784,g2579);
  NR4 NOR4_34(g9876,g9522,g9536,g9576,I15039);
  NR4 NOR4_35(g9656,g9010,g9240,g9223,I14779);
  NR2 NOR2_84(g8303,g8209,g4811);
  NR2 NOR2_85(g10429,g10326,g3507);
  NR2 NOR2_86(g10428,g10335,g4620);
  NR4 NOR4_36(g4234,g3292,g3793,g2586,g3776);
  NR4 NOR4_37(g9877,g9512,g9536,g9569,I15042);
  NR2 NOR2_87(g5186,g2047,g4401);
  NR2 NOR2_88(g9489,g9052,g9030);
  NR4 NOR4_38(g4619,g3077,g3491,g3485,g2655);
  NR2 NOR2_89(g10432,g10350,g3566);
  NR2 NOR2_90(g5345,g2754,g4835);
  NR2 NOR2_91(g5763,g5350,g5345);
  NR2 NOR2_92(g10375,g10288,g3463);
  NR4 NOR4_39(g4879,g3292,g2593,g3784,g2579);
  NR4 NOR4_40(g4607,g3077,g2669,g3485,g3479);
  NR2 NOR2_93(g10425,g10293,g4620);
  NR2 NOR2_94(g3107,g2501,g2499);
  NR2 NOR2_95(g10322,g9317,g10272);
  NR4 NOR4_41(g4630,g3077,g3491,g3485,g3479);
  NR2 NOR2_96(g10364,g10327,g3744);
  NR2 NOR2_97(g9781,g9392,g9367);

endmodule
