module s1196(VDD,CK,G0,G1,G10,G11,G12,G13,G2,G3,G4,G45,G5,G530,G532,G535,
  G537,G539,
  G542,G546,G547,G548,G549,G550,G551,G552,G6,G7,G8,G9);
input VDD,CK,G0,G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13;
output G546,G539,G550,G551,G552,G547,G548,G549,G530,G45,G542,G532,G535,G537;

  wire G29,G502,G30,G503,G31,G504,G32,G505,G33,G506,G34,G507,G35,G508,G36,G509,
    G37,G510,G38,G511,G39,G512,G40,G513,G41,G514,G42,G515,G43,G516,G44,G517,
    G518,G46,G519,G520,G521,G522,G524,II156,G334,G527,G528,G529,G531,G533,G536,
    G538,G540,G541,G543,G476,G484,G125,G140,G132,G70,G67,G99,G475,G57,G59,G58,
    G228,G272,G271,G98,G97,G135,G134,II218,G333,G55,G54,G165,G72,G71,G236,G274,
    G275,II249,G370,G75,G74,G490,G190,G482,G241,G153,G192,G193,G123,G122,II272,
    G209,G458,II276,G238,G332,II280,G309,II287,G347,G498,G195,G78,G77,II295,
    G198,G459,G199,G200,G90,G89,G221,G222,G223,G224,II316,G239,G369,G234,G235,
    II327,G435,II330,G441,G50,G49,G130,G501,G156,G477,G276,G485,II352,G299,
    G497,G205,II371,G335,II374,G456,G87,G86,II386,G414,G486,G68,G231,G232,G160,
    G161,G265,G64,G63,G180,G181,G107,G207,G208,G167,G168,G124,G206,G203,G204,
    G489,G273,G495,G177,G357,G212,G213,II493,G218,G404,II502,G468,G173,G487,
    G534,II529,G149,II536,G79,G446,G494,G500,G214,G215,G492,G62,G483,G182,G282,
    G281,II573,G176,G403,II576,G175,G447,G479,G194,G491,G554,G553,G170,G171,
    G172,G525,G526,G493,G544,G545,G488,G499,G280,II624,G120,G303,G480,G179,
    II631,G188,G336,G496,G174,II662,G405,G478,G279,II692,G145,G432,G359,G469,
    G163,G461,G431,G362,G129,G81,G288,G240,G348,G352,G164,G379,G211,G385,G376,
    G387,G462,G436,G363,G410,G399,G437,G66,G229,G307,G104,G306,G283,G219,G339,
    G472,G136,G351,G169,G440,G382,G100,G386,G85,G321,G378,G471,G191,G103,G112,
    G377,G56,G358,G83,G400,G277,G308,G151,G411,G48,G413,G197,G201,G434,G373,
    G444,G361,G202,G346,G82,G457,G364,G109,G445,G53,G225,G412,G371,G267,G353,
    G92,G388,G114,G473,G143,G331,G257,G429,G51,G380,G93,G360,G106,G338,G337,
    G270,G340,G322,G105,G196,G330,G248,G249,G430,G344,G111,G189,G428,G227,G349,
    G108,G460,G115,G463,G148,G393,G127,G470,G341,G118,G342,G73,G324,G183,G323,
    G144,G354,G312,G315,G250,G251,G474,G242,G343,G147,G304,G52,G158,G398,G94,
    G365,G137,G417,G290,G117,G157,G327,G367,G126,G397,G101,G451,G187,G406,G418,
    G60,G453,G186,G289,G119,G311,G178,G402,G154,G433,G91,G449,G88,G452,G184,
    G329,G150,G291,G138,G155,G328,G102,G366,G372,G116,G383,G131,G392,G396,G76,
    G401,G110,G422,G80,G415,G146,G142,G425,G438,G133,G424,G439,G317,G159,G245,
    G426,G162,G443,G47,G416,G61,G427,G95,G442,G121,G423,G128,G448,G139,G419,
    G394,G407,G314,G395,G302,G355,G316,G350,G368,G381,G384,G389,G374,G286,G293,
    G375,G356,G313,G420,G421,G320,G310,G408,G305,G409,G296,G325,G464,G391,G220,
    G292,G345,G226,G465,G210,G454,G269,G287,G318,G326,G390,G298,G300,G261,G301,
    G297,G455,G152,G319,G284,G294,G141,G285,G295,G450,G244,G166,G252,G216,G263,
    G233,G243,G237,G96,G278,G255,G69,G264,G84,G258,G259,G217,G230,G260,G266,
    G262,G256,G113,G268,G253,G254,G523,G247,G246,G185;

  FD1 DFF_0(CK,G29,G502);
  FD1 DFF_1(CK,G30,G503);
  FD1 DFF_2(CK,G31,G504);
  FD1 DFF_3(CK,G32,G505);
  FD1 DFF_4(CK,G33,G506);
  FD1 DFF_5(CK,G34,G507);
  FD1 DFF_6(CK,G35,G508);
  FD1 DFF_7(CK,G36,G509);
  FD1 DFF_8(CK,G37,G510);
  FD1 DFF_9(CK,G38,G511);
  FD1 DFF_10(CK,G39,G512);
  FD1 DFF_11(CK,G40,G513);
  FD1 DFF_12(CK,G41,G514);
  FD1 DFF_13(CK,G42,G515);
  FD1 DFF_14(CK,G43,G516);
  FD1 DFF_15(CK,G44,G517);
  FD1 DFF_16(CK,G45,G518);
  FD1 DFF_17(CK,G46,G519);
  IV  NOT_0(G520,G0);
  IV  NOT_1(G521,G1);
  IV  NOT_2(G522,G2);
  IV  NOT_3(G524,G3);
  IV  NOT_4(II156,G4);
  IV  NOT_5(G334,II156);
  IV  NOT_6(G527,G4);
  IV  NOT_7(G528,G5);
  IV  NOT_8(G529,G6);
  IV  NOT_9(G531,G7);
  IV  NOT_10(G533,G8);
  IV  NOT_11(G536,G9);
  IV  NOT_12(G538,G10);
  IV  NOT_13(G540,G11);
  IV  NOT_14(G541,G12);
  IV  NOT_15(G543,G13);
  IV  NOT_16(G476,G30);
  IV  NOT_17(G484,G30);
  IV  NOT_18(G125,G40);
  IV  NOT_19(G140,G33);
  IV  NOT_20(G546,G41);
  IV  NOT_21(G132,G42);
  IV  NOT_22(G70,G43);
  IV  NOT_23(G67,G44);
  IV  NOT_24(G99,G29);
  IV  NOT_25(G475,G57);
  IV  NOT_26(G59,G58);
  IV  NOT_27(G228,G524);
  IV  NOT_28(G272,G271);
  IV  NOT_29(G98,G97);
  IV  NOT_30(G135,G134);
  IV  NOT_31(II218,G528);
  IV  NOT_32(G333,II218);
  IV  NOT_33(G55,G54);
  IV  NOT_34(G165,G529);
  IV  NOT_35(G72,G71);
  IV  NOT_36(G236,G274);
  IV  NOT_37(G275,G274);
  IV  NOT_38(II249,G538);
  IV  NOT_39(G370,II249);
  IV  NOT_40(G75,G74);
  IV  NOT_41(G490,G190);
  IV  NOT_42(G482,G241);
  IV  NOT_43(G153,G522);
  IV  NOT_44(G192,G193);
  IV  NOT_45(G123,G122);
  IV  NOT_46(II272,G209);
  IV  NOT_47(G458,II272);
  IV  NOT_48(II276,G238);
  IV  NOT_49(G332,II276);
  IV  NOT_50(II280,G272);
  IV  NOT_51(G309,II280);
  IV  NOT_52(II287,G135);
  IV  NOT_53(G347,II287);
  IV  NOT_54(G498,G195);
  IV  NOT_55(G78,G77);
  IV  NOT_56(II295,G198);
  IV  NOT_57(G459,II295);
  IV  NOT_58(G199,G200);
  IV  NOT_59(G90,G89);
  IV  NOT_60(G221,G222);
  IV  NOT_61(G223,G224);
  IV  NOT_62(II316,G239);
  IV  NOT_63(G369,II316);
  IV  NOT_64(G234,G235);
  IV  NOT_65(II327,G135);
  IV  NOT_66(G435,II327);
  IV  NOT_67(II330,G236);
  IV  NOT_68(G441,II330);
  IV  NOT_69(G50,G49);
  IV  NOT_70(G130,G9);
  IV  NOT_71(G501,G156);
  IV  NOT_72(G477,G276);
  IV  NOT_73(G485,G276);
  IV  NOT_74(II352,G77);
  IV  NOT_75(G299,II352);
  IV  NOT_76(G497,G205);
  IV  NOT_77(II371,G1);
  IV  NOT_78(G335,II371);
  IV  NOT_79(II374,G520);
  IV  NOT_80(G456,II374);
  IV  NOT_81(G87,G86);
  IV  NOT_82(II386,G199);
  IV  NOT_83(G414,II386);
  IV  NOT_84(G486,G68);
  IV  NOT_85(G231,G232);
  IV  NOT_86(G160,G161);
  IV  NOT_87(G265,G50);
  IV  NOT_88(G64,G63);
  IV  NOT_89(G180,G181);
  IV  NOT_90(G107,G456);
  IV  NOT_91(G207,G208);
  IV  NOT_92(G167,G168);
  IV  NOT_93(G124,G206);
  IV  NOT_94(G203,G204);
  IV  NOT_95(G489,G273);
  IV  NOT_96(G495,G273);
  IV  NOT_97(G177,G357);
  IV  NOT_98(G212,G213);
  IV  NOT_99(II493,G218);
  IV  NOT_100(G404,II493);
  IV  NOT_101(II502,G124);
  IV  NOT_102(G468,II502);
  IV  NOT_103(G173,G495);
  IV  NOT_104(G487,G534);
  IV  NOT_105(II529,G468);
  IV  NOT_106(G149,II529);
  IV  NOT_107(II536,G79);
  IV  NOT_108(G446,II536);
  IV  NOT_109(G494,G173);
  IV  NOT_110(G500,G173);
  IV  NOT_111(G214,G215);
  IV  NOT_112(G492,G62);
  IV  NOT_113(G483,G182);
  IV  NOT_114(G282,G281);
  IV  NOT_115(II573,G176);
  IV  NOT_116(G403,II573);
  IV  NOT_117(II576,G175);
  IV  NOT_118(G447,II576);
  IV  NOT_119(G479,G194);
  IV  NOT_120(G491,G194);
  IV  NOT_121(G554,G553);
  IV  NOT_122(G170,G171);
  IV  NOT_123(G172,G171);
  IV  NOT_124(G525,G526);
  IV  NOT_125(G493,G544);
  IV  NOT_126(G545,G544);
  IV  NOT_127(G488,G172);
  IV  NOT_128(G499,G280);
  IV  NOT_129(II624,G120);
  IV  NOT_130(G303,II624);
  IV  NOT_131(G480,G179);
  IV  NOT_132(II631,G188);
  IV  NOT_133(G336,II631);
  IV  NOT_134(G496,G188);
  IV  NOT_135(G174,G496);
  IV  NOT_136(II662,G174);
  IV  NOT_137(G405,II662);
  IV  NOT_138(G478,G279);
  IV  NOT_139(II692,G145);
  IV  NOT_140(G432,II692);
  AN2 AND2_0(G359,G6,G31);
  AN2 AND2_1(G469,G163,G3);
  AN2 AND2_2(G461,G529,G531);
  AN2 AND2_3(G431,G524,G67);
  AN2 AND2_4(G362,G129,G77);
  AN2 AND2_5(G81,G288,G240);
  AN2 AND2_6(G348,G97,G55);
  AN4 AND4_0(G352,G8,G135,G37,G164);
  AN2 AND2_7(G511,G163,G164);
  AN2 AND2_8(G379,G9,G211);
  AN3 AND3_0(G385,G529,G7,G49);
  AN2 AND2_9(G376,G533,G75);
  AN3 AND3_1(G387,G6,G274,G75);
  AN2 AND2_10(G462,G192,G538);
  AN2 AND2_11(G436,G123,G77);
  AN2 AND2_12(G363,G77,G205);
  AN2 AND2_13(G410,G1,G205);
  AN2 AND2_14(G399,G520,G1);
  AN2 AND2_15(G437,G66,G229);
  AN2 AND2_16(G307,G6,G104);
  AN2 AND2_17(G306,G524,G78);
  AN2 AND2_18(G283,G122,G219);
  AN3 AND3_2(G339,G533,G199,G209);
  AN3 AND3_3(G472,G136,G9,G190);
  AN4 AND4_1(G351,G524,G169,G221,G234);
  AN2 AND2_19(G440,G38,G234);
  AN3 AND3_4(G382,G9,G100,G34);
  AN2 AND2_20(G386,G536,G85);
  AN2 AND2_21(G321,G90,G50);
  AN2 AND2_22(G378,G89,G50);
  AN3 AND3_5(G471,G191,G103,G112);
  AN2 AND2_23(G377,G90,G56);
  AN2 AND2_24(G358,G7,G83);
  AN2 AND2_25(G400,G0,G277);
  AN2 AND2_26(G308,G5,G151);
  AN2 AND2_27(G411,G48,G59);
  AN2 AND2_28(G413,G197,G201);
  AN2 AND2_29(G434,G165,G231);
  AN2 AND2_30(G373,G34,G160);
  AN2 AND2_31(G357,G265,G232);
  AN3 AND3_6(G444,G64,G78,G211);
  AN2 AND2_32(G361,G6,G202);
  AN2 AND2_33(G346,G2,G82);
  AN2 AND2_34(G457,G4,G107);
  AN2 AND2_35(G364,G2,G109);
  AN2 AND2_36(G445,G53,G225);
  AN2 AND2_37(G412,G3,G207);
  AN3 AND3_7(G371,G161,G168,G267);
  AN3 AND3_8(G353,G11,G92,G163);
  AN2 AND2_38(G388,G11,G114);
  AN2 AND2_39(G473,G11,G143);
  AN2 AND2_40(G331,G213,G257);
  AN2 AND2_41(G429,G51,G225);
  AN2 AND2_42(G380,G6,G93);
  AN2 AND2_43(G360,G8,G106);
  AN2 AND2_44(G338,G202,G203);
  AN2 AND2_45(G337,G270,G167);
  AN2 AND2_46(G340,G8,G270);
  AN3 AND3_9(G322,G522,G105,G196);
  AN2 AND2_47(G330,G248,G249);
  AN2 AND2_48(G430,G177,G196);
  AN3 AND3_10(G344,G111,G189,G195);
  AN2 AND2_49(G428,G212,G227);
  AN2 AND2_50(G349,G6,G108);
  AN3 AND3_11(G460,G2,G81,G115);
  AN2 AND2_51(G463,G521,G148);
  AN2 AND2_52(G393,G127,G34);
  AN2 AND2_53(G470,G528,G149);
  AN2 AND2_54(G341,G531,G118);
  AN2 AND2_55(G342,G73,G197);
  AN2 AND2_56(G324,G522,G183);
  AN2 AND2_57(G323,G2,G144);
  AN2 AND2_58(G354,G0,G214);
  AN2 AND2_59(G312,G180,G182);
  AN2 AND2_60(G315,G250,G251);
  AN2 AND2_61(G474,G242,G77);
  AN3 AND3_12(G343,G2,G528,G147);
  AN2 AND2_62(G304,G52,G158);
  AN3 AND3_13(G398,G94,G156,G158);
  AN3 AND3_14(G365,G282,G137,G156);
  AN3 AND3_15(G417,G13,G282,G70);
  AN3 AND3_16(G290,G117,G135,G157);
  AN3 AND3_17(G327,G4,G39,G157);
  AN2 AND2_63(G367,G126,G157);
  AN3 AND3_18(G397,G101,G98,G157);
  AN3 AND3_19(G451,G541,G554,G187);
  AN2 AND2_64(G406,G87,G172);
  AN3 AND3_20(G418,G524,G60,G172);
  AN2 AND2_65(G453,G545,G186);
  AN3 AND3_21(G289,G2,G119,G156);
  AN3 AND3_22(G311,G0,G178,G179);
  AN2 AND2_66(G402,G154,G183);
  AN2 AND2_67(G433,G91,G154);
  AN2 AND2_68(G449,G88,G154);
  AN2 AND2_69(G452,G526,G184);
  AN2 AND2_70(G329,G150,G156);
  AN2 AND2_71(G291,G138,G155);
  AN3 AND3_23(G328,G5,G102,G155);
  AN2 AND2_72(G366,G125,G155);
  AN3 AND3_24(G372,G116,G275,G155);
  AN2 AND2_73(G383,G131,G155);
  AN2 AND2_74(G392,G132,G155);
  AN3 AND3_25(G396,G76,G272,G155);
  AN3 AND3_26(G401,G2,G110,G155);
  AN3 AND3_27(G422,G0,G80,G155);
  AN3 AND3_28(G415,G146,G142,G165);
  AN2 AND2_75(G425,G146,G176);
  AN3 AND3_29(G438,G8,G146,G133);
  AN3 AND3_30(G424,G78,G174,G177);
  AN2 AND2_76(G439,G174,G175);
  AN2 AND2_77(G317,G159,G245);
  AN3 AND3_31(G426,G37,G162,G38);
  AN2 AND2_78(G443,G47,G162);
  AN2 AND2_79(G416,G61,G167);
  AN3 AND3_32(G427,G541,G95,G165);
  AN2 AND2_80(G442,G541,G121);
  AN2 AND2_81(G423,G541,G128);
  AN2 AND2_82(G448,G139,G153);
  OR2 OR2_0(G419,G3,G5);
  OR2 OR2_1(G193,G6,G30);
  OR2 OR2_2(G394,G5,G58);
  OR2 OR2_3(G407,G6,G117);
  OR2 OR2_4(G314,G527,G57);
  OR2 OR2_5(G395,G4,G134);
  OR2 OR2_6(G288,G1,G528);
  OR2 OR2_7(G302,G4,G529);
  OR2 OR2_8(G224,G533,G31);
  OR2 OR2_9(G355,G11,G116);
  OR2 OR2_10(G316,G531,G536);
  OR2 OR2_11(G350,G6,G536);
  OR2 OR2_12(G368,G533,G536);
  OR2 OR2_13(G381,G7,G71);
  OR2 OR2_14(G384,G529,G71);
  OR2 OR2_15(G389,G9,G274);
  OR2 OR2_16(G374,G536,G538);
  OR2 OR2_17(G286,G9,G540);
  OR2 OR2_18(G293,G7,G540);
  OR2 OR2_19(G375,G10,G540);
  OR2 OR2_20(G356,G6,G476);
  OR2 OR2_21(G313,G521,G475);
  OR2 OR2_22(G420,G522,G59);
  OR3 OR3_0(G421,G521,G2,G228);
  OR2 OR2_23(G320,G76,G272);
  OR2 OR2_24(G310,G522,G135);
  OR2 OR2_25(G408,G529,G77);
  OR2 OR2_26(G305,G524,G55);
  OR2 OR2_27(G409,G528,G55);
  OR2 OR2_28(G296,G89,G484);
  OR3 OR3_1(G325,G7,G536,G222);
  OR2 OR2_29(G464,G72,G536);
  OR2 OR2_30(G391,G74,G220);
  OR2 OR2_31(G292,G538,G75);
  OR2 OR2_32(G345,G529,G226);
  OR2 OR2_33(G465,G524,G210);
  OR2 OR2_34(G454,G122,G77);
  OR2 OR2_35(G269,G362,G529);
  OR2 OR2_36(G287,G522,G81);
  OR3 OR3_2(G318,G6,G8,G232);
  OR2 OR2_37(G326,G533,G232);
  OR2 OR2_38(G390,G89,G50);
  OR2 OR2_39(G298,G5,G497);
  OR2 OR2_40(G300,G87,G97);
  OR2 OR2_41(G261,G283,G528);
  OR2 OR2_42(G301,G122,G486);
  OR2 OR2_43(G92,G351,G352);
  OR2 OR2_44(G47,G440,G441);
  OR2 OR2_45(G114,G385,G386);
  OR2 OR2_46(G297,G64,G274);
  OR3 OR3_3(G93,G376,G377,G378);
  OR2 OR2_47(G106,G358,G359);
  OR2 OR2_48(G110,G399,G400);
  OR2 OR2_49(G455,G78,G206);
  OR3 OR3_4(G152,G306,G307,G308);
  OR2 OR2_50(G60,G413,G414);
  OR2 OR2_51(G133,G434,G435);
  OR2 OR2_52(G105,G321,G273);
  OR2 OR2_53(G108,G346,G347);
  OR3 OR3_5(G115,G457,G458,G459);
  OR2 OR2_54(G126,G363,G364);
  OR2 OR2_55(G79,G444,G445);
  OR2 OR2_56(G319,G529,G489);
  OR2 OR2_57(G131,G379,G380);
  OR2 OR2_58(G118,G337,G338);
  OR2 OR2_59(G73,G339,G340);
  OR2 OR2_60(G91,G430,G431);
  OR2 OR2_61(G137,G348,G349);
  OR2 OR2_62(G242,G469,G470);
  OR2 OR2_63(G147,G341,G342);
  OR3 OR3_6(G284,G528,G272,G281);
  OR3 OR3_7(G294,G1,G117,G281);
  OR3 OR3_8(G553,G322,G323,G324);
  OR2 OR2_64(G141,G353,G354);
  OR2 OR2_65(G142,G403,G404);
  OR2 OR2_66(G88,G446,G447);
  OR2 OR2_67(G544,G343,G344);
  OR2 OR2_68(G285,G5,G479);
  OR2 OR2_69(G295,G122,G491);
  OR2 OR2_70(G450,G12,G171);
  OR2 OR2_71(G150,G303,G304);
  OR2 OR2_72(G146,G336,G170);
  OR3 OR3_9(G539,G451,G452,G453);
  OR2 OR2_73(G244,G371,G159);
  OR4 OR4_0(G550,G289,G290,G291,G485);
  OR3 OR3_10(G551,G327,G328,G329);
  OR3 OR3_11(G552,G365,G366,G367);
  OR2 OR2_74(G547,G382,G383);
  OR2 OR2_75(G548,G392,G393);
  OR4 OR4_1(G549,G396,G397,G398,G477);
  OR2 OR2_76(G530,G401,G402);
  OR2 OR2_77(G61,G405,G406);
  OR2 OR2_78(G95,G424,G425);
  OR2 OR2_79(G121,G438,G439);
  OR2 OR2_80(G279,G317,G166);
  OR4 OR4_2(G128,G415,G416,G417,G418);
  OR2 OR2_81(G145,G426,G427);
  OR2 OR2_82(G139,G442,G443);
  OR2 OR2_83(G532,G422,G423);
  OR2 OR2_84(G535,G432,G433);
  OR2 OR2_85(G537,G448,G449);
  ND2 NAND2_0(G57,G0,G2);
  ND2 NAND2_1(G58,G1,G3);
  ND2 NAND2_2(G76,G0,G3);
  ND2 NAND2_3(G101,G3,G4);
  ND2 NAND2_4(G117,G2,G4);
  ND2 NAND2_5(G271,G1,G4);
  ND2 NAND2_6(G97,G2,G5);
  ND2 NAND2_7(G134,G3,G5);
  ND2 NAND2_8(G54,G4,G6);
  ND2 NAND2_9(G116,G6,G9);
  ND2 NAND2_10(G71,G8,G10);
  ND2 NAND2_11(G274,G7,G10);
  ND2 NAND2_12(G74,G9,G11);
  ND2 NAND2_13(G112,G8,G31);
  ND2 NAND2_14(G245,G8,G34);
  ND2 NAND2_15(G122,G522,G3);
  ND2 NAND2_16(G238,G2,G524);
  ND2 NAND2_17(G129,G527,G5);
  ND2 NAND2_18(G240,G4,G134);
  ND4 NAND4_0(G252,G3,G11,G35,G216);
  ND2 NAND2_19(G77,G4,G528);
  ND3 NAND3_0(G103,G529,G7,G30);
  ND2 NAND2_20(G200,G527,G529);
  ND2 NAND2_21(G248,G529,G36);
  ND2 NAND2_22(G89,G531,G8);
  ND2 NAND2_23(G222,G533,G10);
  ND2 NAND2_24(G239,G7,G533);
  ND2 NAND2_25(G235,G6,G536);
  ND2 NAND2_26(G220,G7,G71);
  ND2 NAND2_27(G49,G9,G538);
  ND2 NAND2_28(G251,G543,G32);
  ND3 NAND3_1(G276,G3,G543,G140);
  ND2 NAND2_29(G263,G0,G99);
  ND2 NAND2_30(G226,G527,G59);
  ND2 NAND2_31(G210,G520,G272);
  ND2 NAND2_32(G66,G129,G101);
  ND2 NAND2_33(G233,G522,G135);
  ND3 NAND3_2(G104,G122,G238,G240);
  ND2 NAND2_34(G86,G55,G3);
  ND2 NAND2_35(G219,G524,G55);
  ND2 NAND2_36(G68,G302,G528);
  ND2 NAND2_37(G232,G536,G164);
  ND2 NAND2_38(G136,G222,G224);
  ND2 NAND2_39(G510,G350,G235);
  ND2 NAND2_40(G161,G316,G72);
  ND2 NAND2_41(G100,G381,G220);
  ND2 NAND2_42(G85,G384,G239);
  ND3 NAND3_3(G243,G368,G275,G34);
  ND2 NAND2_43(G63,G75,G8);
  ND3 NAND3_4(G237,G10,G75,G201);
  ND2 NAND2_44(G503,G286,G538);
  ND2 NAND2_45(G56,G374,G375);
  ND2 NAND2_46(G83,G355,G356);
  ND2 NAND2_47(G96,G313,G314);
  ND2 NAND2_48(G278,G332,G333);
  ND3 NAND3_5(G255,G309,G2,G529);
  ND3 NAND3_6(G69,G419,G420,G233);
  ND2 NAND2_49(G512,G310,G233);
  ND2 NAND2_50(G181,G2,G78);
  ND3 NAND3_7(G277,G394,G395,G81);
  ND2 NAND2_51(G151,G305,G200);
  ND3 NAND3_8(G48,G407,G408,G409);
  ND2 NAND2_52(G264,G227,G241);
  ND2 NAND2_53(G208,G68,G229);
  ND2 NAND2_54(G168,G75,G221);
  ND2 NAND2_55(G84,G369,G370);
  ND3 NAND3_9(G258,G464,G103,G223);
  ND2 NAND2_56(G166,G7,G50);
  ND2 NAND2_57(G259,G130,G225);
  ND2 NAND2_58(G504,G292,G293);
  ND2 NAND2_59(G217,G50,G230);
  ND2 NAND2_60(G257,G538,G230);
  ND3 NAND3_10(G260,G528,G529,G191);
  ND2 NAND2_61(G266,G524,G96);
  ND2 NAND2_62(G262,G527,G278);
  ND2 NAND2_63(G138,G465,G263);
  ND2 NAND2_64(G256,G4,G69);
  ND2 NAND2_65(G82,G334,G335);
  ND2 NAND2_66(G109,G269,G219);
  ND2 NAND2_67(G206,G287,G524);
  ND2 NAND2_68(G204,G521,G87);
  ND2 NAND2_69(G53,G264,G237);
  ND2 NAND2_70(G273,G325,G326);
  ND2 NAND2_71(G267,G536,G84);
  ND2 NAND2_72(G113,G389,G390);
  ND3 NAND3_11(G143,G258,G193,G259);
  ND2 NAND2_73(G213,G64,G275);
  ND2 NAND2_74(G51,G260,G237);
  ND3 NAND3_12(G102,G320,G266,G210);
  ND3 NAND3_13(G52,G298,G299,G219);
  ND3 NAND3_14(G80,G421,G226,G256);
  ND2 NAND2_75(G270,G345,G204);
  ND3 NAND3_15(G94,G261,G181,G262);
  ND3 NAND3_16(G505,G300,G301,G181);
  ND3 NAND3_17(G249,G11,G273,G201);
  ND2 NAND2_76(G268,G11,G113);
  ND2 NAND2_77(G111,G213,G217);
  ND3 NAND3_18(G534,G296,G297,G166);
  ND2 NAND2_78(G253,G87,G218);
  ND3 NAND3_19(G148,G454,G455,G0);
  ND2 NAND2_79(G254,G1,G152);
  ND2 NAND2_80(G127,G391,G268);
  ND3 NAND3_20(G215,G135,G55,G212);
  ND2 NAND2_81(G62,G534,G32);
  ND3 NAND3_21(G523,G254,G255,G208);
  ND2 NAND2_82(G508,G318,G319);
  ND3 NAND3_22(G144,G215,G252,G253);
  ND2 NAND2_83(G250,G13,G523);
  ND2 NAND2_84(G281,G523,G534);
  ND2 NAND2_85(G171,G553,G187);
  ND3 NAND3_23(G526,G1,G2,G141);
  ND2 NAND2_86(G280,G46,G247);
  ND2 NAND2_87(G246,G544,G186);
  ND2 NAND2_88(G119,G284,G285);
  ND2 NAND2_89(G120,G294,G295);
  ND2 NAND2_90(G185,G525,G184);
  ND2 NAND2_91(G159,G6,G155);
  ND3 NAND3_24(G518,G450,G185,G246);
  ND3 NAND3_25(G542,G243,G244,G279);
  NR2 NOR2_0(G163,G0,G4);
  NR2 NOR2_1(G216,G4,G5);
  NR2 NOR2_2(G169,G5,G7);
  NR2 NOR2_3(G225,G7,G8);
  NR2 NOR2_4(G190,G7,G11);
  NR2 NOR2_5(G241,G10,G11);
  NR2 NOR2_6(G198,G520,G3);
  NR2 NOR2_7(G178,G521,G4);
  NR2 NOR2_8(G229,G1,G522);
  NR2 NOR2_9(G209,G1,G524);
  NR2 NOR2_10(G195,G521,G134);
  NR2 NOR2_11(G189,G522,G54);
  NR2 NOR2_12(G201,G528,G54);
  NR2 NOR2_13(G164,G531,G10);
  NR2 NOR2_14(G211,G6,G274);
  NR2 NOR2_15(G156,G12,G543);
  NR2 NOR2_16(G205,G529,G122);
  NR2 NOR2_17(G227,G5,G200);
  NR2 NOR2_18(G230,G8,G490);
  NR2 NOR2_19(G191,G9,G482);
  NR3 NOR3_0(G196,G5,G540,G86);
  NR2 NOR2_20(G197,G540,G232);
  NR2 NOR2_21(G202,G10,G63);
  NR2 NOR2_22(G502,G436,G437);
  NR2 NOR2_23(G218,G528,G217);
  NR3 NOR3_1(G516,G410,G411,G412);
  NR2 NOR2_24(G515,G387,G388);
  NR2 NOR2_25(G509,G331,G5);
  NR2 NOR2_26(G513,G360,G361);
  NR2 NOR2_27(G183,G330,G3);
  NR2 NOR2_28(G517,G428,G429);
  NR2 NOR2_29(G182,G12,G62);
  NR4 NOR4_0(G519,G460,G461,G462,G463);
  NR2 NOR2_30(G176,G4,G494);
  NR2 NOR2_31(G175,G86,G500);
  NR2 NOR2_32(G187,G13,G492);
  NR2 NOR2_33(G158,G521,G281);
  NR2 NOR2_34(G194,G281,G271);
  NR2 NOR2_35(G157,G13,G483);
  NR3 NOR3_2(G507,G315,G12,G487);
  NR2 NOR2_36(G186,G282,G501);
  NR4 NOR4_1(G247,G471,G472,G473,G474);
  NR2 NOR2_37(G179,G541,G280);
  NR2 NOR2_38(G188,G543,G493);
  NR2 NOR2_39(G154,G12,G488);
  NR3 NOR3_3(G184,G541,G13,G499);
  NR2 NOR2_40(G506,G311,G312);
  NR2 NOR2_41(G155,G13,G480);
  NR2 NOR2_42(G162,G185,G498);
  NR3 NOR3_4(G514,G372,G373,G478);

endmodule
